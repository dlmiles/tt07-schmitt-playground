magic
tech sky130A
magscale 1 2
timestamp 1716692466
<< error_p >>
rect -287 472 -225 478
rect -159 472 -97 478
rect -31 472 31 478
rect 97 472 159 478
rect 225 472 287 478
rect -287 438 -275 472
rect -159 438 -147 472
rect -31 438 -19 472
rect 97 438 109 472
rect 225 438 237 472
rect -287 432 -225 438
rect -159 432 -97 438
rect -31 432 31 438
rect 97 432 159 438
rect 225 432 287 438
rect -287 -438 -225 -432
rect -159 -438 -97 -432
rect -31 -438 31 -432
rect 97 -438 159 -432
rect 225 -438 287 -432
rect -287 -472 -275 -438
rect -159 -472 -147 -438
rect -31 -472 -19 -438
rect 97 -472 109 -438
rect 225 -472 237 -438
rect -287 -478 -225 -472
rect -159 -478 -97 -472
rect -31 -478 31 -472
rect 97 -478 159 -472
rect 225 -478 287 -472
<< pwell >>
rect -487 -610 487 610
<< nmoslvt >>
rect -291 -400 -221 400
rect -163 -400 -93 400
rect -35 -400 35 400
rect 93 -400 163 400
rect 221 -400 291 400
<< ndiff >>
rect -349 388 -291 400
rect -349 -388 -337 388
rect -303 -388 -291 388
rect -349 -400 -291 -388
rect -221 388 -163 400
rect -221 -388 -209 388
rect -175 -388 -163 388
rect -221 -400 -163 -388
rect -93 388 -35 400
rect -93 -388 -81 388
rect -47 -388 -35 388
rect -93 -400 -35 -388
rect 35 388 93 400
rect 35 -388 47 388
rect 81 -388 93 388
rect 35 -400 93 -388
rect 163 388 221 400
rect 163 -388 175 388
rect 209 -388 221 388
rect 163 -400 221 -388
rect 291 388 349 400
rect 291 -388 303 388
rect 337 -388 349 388
rect 291 -400 349 -388
<< ndiffc >>
rect -337 -388 -303 388
rect -209 -388 -175 388
rect -81 -388 -47 388
rect 47 -388 81 388
rect 175 -388 209 388
rect 303 -388 337 388
<< psubdiff >>
rect -451 540 -355 574
rect 355 540 451 574
rect -451 478 -417 540
rect 417 478 451 540
rect -451 -540 -417 -478
rect 417 -540 451 -478
rect -451 -574 -355 -540
rect 355 -574 451 -540
<< psubdiffcont >>
rect -355 540 355 574
rect -451 -478 -417 478
rect 417 -478 451 478
rect -355 -574 355 -540
<< poly >>
rect -291 472 -221 488
rect -291 438 -275 472
rect -237 438 -221 472
rect -291 400 -221 438
rect -163 472 -93 488
rect -163 438 -147 472
rect -109 438 -93 472
rect -163 400 -93 438
rect -35 472 35 488
rect -35 438 -19 472
rect 19 438 35 472
rect -35 400 35 438
rect 93 472 163 488
rect 93 438 109 472
rect 147 438 163 472
rect 93 400 163 438
rect 221 472 291 488
rect 221 438 237 472
rect 275 438 291 472
rect 221 400 291 438
rect -291 -438 -221 -400
rect -291 -472 -275 -438
rect -237 -472 -221 -438
rect -291 -488 -221 -472
rect -163 -438 -93 -400
rect -163 -472 -147 -438
rect -109 -472 -93 -438
rect -163 -488 -93 -472
rect -35 -438 35 -400
rect -35 -472 -19 -438
rect 19 -472 35 -438
rect -35 -488 35 -472
rect 93 -438 163 -400
rect 93 -472 109 -438
rect 147 -472 163 -438
rect 93 -488 163 -472
rect 221 -438 291 -400
rect 221 -472 237 -438
rect 275 -472 291 -438
rect 221 -488 291 -472
<< polycont >>
rect -275 438 -237 472
rect -147 438 -109 472
rect -19 438 19 472
rect 109 438 147 472
rect 237 438 275 472
rect -275 -472 -237 -438
rect -147 -472 -109 -438
rect -19 -472 19 -438
rect 109 -472 147 -438
rect 237 -472 275 -438
<< locali >>
rect -451 540 -355 574
rect 355 540 451 574
rect -451 478 -417 540
rect 417 478 451 540
rect -291 438 -275 472
rect -237 438 -221 472
rect -163 438 -147 472
rect -109 438 -93 472
rect -35 438 -19 472
rect 19 438 35 472
rect 93 438 109 472
rect 147 438 163 472
rect 221 438 237 472
rect 275 438 291 472
rect -337 388 -303 404
rect -337 -404 -303 -388
rect -209 388 -175 404
rect -209 -404 -175 -388
rect -81 388 -47 404
rect -81 -404 -47 -388
rect 47 388 81 404
rect 47 -404 81 -388
rect 175 388 209 404
rect 175 -404 209 -388
rect 303 388 337 404
rect 303 -404 337 -388
rect -291 -472 -275 -438
rect -237 -472 -221 -438
rect -163 -472 -147 -438
rect -109 -472 -93 -438
rect -35 -472 -19 -438
rect 19 -472 35 -438
rect 93 -472 109 -438
rect 147 -472 163 -438
rect 221 -472 237 -438
rect 275 -472 291 -438
rect -451 -540 -417 -478
rect 417 -540 451 -478
rect -451 -574 -355 -540
rect 355 -574 451 -540
<< viali >>
rect -275 438 -237 472
rect -147 438 -109 472
rect -19 438 19 472
rect 109 438 147 472
rect 237 438 275 472
rect -337 -388 -303 388
rect -209 -388 -175 388
rect -81 -388 -47 388
rect 47 -388 81 388
rect 175 -388 209 388
rect 303 -388 337 388
rect -275 -472 -237 -438
rect -147 -472 -109 -438
rect -19 -472 19 -438
rect 109 -472 147 -438
rect 237 -472 275 -438
<< metal1 >>
rect -287 472 -225 478
rect -287 438 -275 472
rect -237 438 -225 472
rect -287 432 -225 438
rect -159 472 -97 478
rect -159 438 -147 472
rect -109 438 -97 472
rect -159 432 -97 438
rect -31 472 31 478
rect -31 438 -19 472
rect 19 438 31 472
rect -31 432 31 438
rect 97 472 159 478
rect 97 438 109 472
rect 147 438 159 472
rect 97 432 159 438
rect 225 472 287 478
rect 225 438 237 472
rect 275 438 287 472
rect 225 432 287 438
rect -343 388 -297 400
rect -343 -388 -337 388
rect -303 -388 -297 388
rect -343 -400 -297 -388
rect -215 388 -169 400
rect -215 -388 -209 388
rect -175 -388 -169 388
rect -215 -400 -169 -388
rect -87 388 -41 400
rect -87 -388 -81 388
rect -47 -388 -41 388
rect -87 -400 -41 -388
rect 41 388 87 400
rect 41 -388 47 388
rect 81 -388 87 388
rect 41 -400 87 -388
rect 169 388 215 400
rect 169 -388 175 388
rect 209 -388 215 388
rect 169 -400 215 -388
rect 297 388 343 400
rect 297 -388 303 388
rect 337 -388 343 388
rect 297 -400 343 -388
rect -287 -438 -225 -432
rect -287 -472 -275 -438
rect -237 -472 -225 -438
rect -287 -478 -225 -472
rect -159 -438 -97 -432
rect -159 -472 -147 -438
rect -109 -472 -97 -438
rect -159 -478 -97 -472
rect -31 -438 31 -432
rect -31 -472 -19 -438
rect 19 -472 31 -438
rect -31 -478 31 -472
rect 97 -438 159 -432
rect 97 -472 109 -438
rect 147 -472 159 -438
rect 97 -478 159 -472
rect 225 -438 287 -432
rect 225 -472 237 -438
rect 275 -472 287 -438
rect 225 -478 287 -472
<< properties >>
string FIXED_BBOX -434 -557 434 557
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4 l 0.350 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
