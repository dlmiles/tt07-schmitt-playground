magic
tech sky130A
magscale 1 2
timestamp 1716692466
<< error_p >>
rect -671 681 -609 687
rect -543 681 -481 687
rect -415 681 -353 687
rect -287 681 -225 687
rect -159 681 -97 687
rect -31 681 31 687
rect 97 681 159 687
rect 225 681 287 687
rect 353 681 415 687
rect 481 681 543 687
rect 609 681 671 687
rect -671 647 -659 681
rect -543 647 -531 681
rect -415 647 -403 681
rect -287 647 -275 681
rect -159 647 -147 681
rect -31 647 -19 681
rect 97 647 109 681
rect 225 647 237 681
rect 353 647 365 681
rect 481 647 493 681
rect 609 647 621 681
rect -671 641 -609 647
rect -543 641 -481 647
rect -415 641 -353 647
rect -287 641 -225 647
rect -159 641 -97 647
rect -31 641 31 647
rect 97 641 159 647
rect 225 641 287 647
rect 353 641 415 647
rect 481 641 543 647
rect 609 641 671 647
rect -671 -647 -609 -641
rect -543 -647 -481 -641
rect -415 -647 -353 -641
rect -287 -647 -225 -641
rect -159 -647 -97 -641
rect -31 -647 31 -641
rect 97 -647 159 -641
rect 225 -647 287 -641
rect 353 -647 415 -641
rect 481 -647 543 -641
rect 609 -647 671 -641
rect -671 -681 -659 -647
rect -543 -681 -531 -647
rect -415 -681 -403 -647
rect -287 -681 -275 -647
rect -159 -681 -147 -647
rect -31 -681 -19 -647
rect 97 -681 109 -647
rect 225 -681 237 -647
rect 353 -681 365 -647
rect 481 -681 493 -647
rect 609 -681 621 -647
rect -671 -687 -609 -681
rect -543 -687 -481 -681
rect -415 -687 -353 -681
rect -287 -687 -225 -681
rect -159 -687 -97 -681
rect -31 -687 31 -681
rect 97 -687 159 -681
rect 225 -687 287 -681
rect 353 -687 415 -681
rect 481 -687 543 -681
rect 609 -687 671 -681
<< nwell >>
rect -871 -819 871 819
<< pmoslvt >>
rect -675 -600 -605 600
rect -547 -600 -477 600
rect -419 -600 -349 600
rect -291 -600 -221 600
rect -163 -600 -93 600
rect -35 -600 35 600
rect 93 -600 163 600
rect 221 -600 291 600
rect 349 -600 419 600
rect 477 -600 547 600
rect 605 -600 675 600
<< pdiff >>
rect -733 588 -675 600
rect -733 -588 -721 588
rect -687 -588 -675 588
rect -733 -600 -675 -588
rect -605 588 -547 600
rect -605 -588 -593 588
rect -559 -588 -547 588
rect -605 -600 -547 -588
rect -477 588 -419 600
rect -477 -588 -465 588
rect -431 -588 -419 588
rect -477 -600 -419 -588
rect -349 588 -291 600
rect -349 -588 -337 588
rect -303 -588 -291 588
rect -349 -600 -291 -588
rect -221 588 -163 600
rect -221 -588 -209 588
rect -175 -588 -163 588
rect -221 -600 -163 -588
rect -93 588 -35 600
rect -93 -588 -81 588
rect -47 -588 -35 588
rect -93 -600 -35 -588
rect 35 588 93 600
rect 35 -588 47 588
rect 81 -588 93 588
rect 35 -600 93 -588
rect 163 588 221 600
rect 163 -588 175 588
rect 209 -588 221 588
rect 163 -600 221 -588
rect 291 588 349 600
rect 291 -588 303 588
rect 337 -588 349 588
rect 291 -600 349 -588
rect 419 588 477 600
rect 419 -588 431 588
rect 465 -588 477 588
rect 419 -600 477 -588
rect 547 588 605 600
rect 547 -588 559 588
rect 593 -588 605 588
rect 547 -600 605 -588
rect 675 588 733 600
rect 675 -588 687 588
rect 721 -588 733 588
rect 675 -600 733 -588
<< pdiffc >>
rect -721 -588 -687 588
rect -593 -588 -559 588
rect -465 -588 -431 588
rect -337 -588 -303 588
rect -209 -588 -175 588
rect -81 -588 -47 588
rect 47 -588 81 588
rect 175 -588 209 588
rect 303 -588 337 588
rect 431 -588 465 588
rect 559 -588 593 588
rect 687 -588 721 588
<< nsubdiff >>
rect -835 749 -739 783
rect 739 749 835 783
rect -835 687 -801 749
rect 801 687 835 749
rect -835 -749 -801 -687
rect 801 -749 835 -687
rect -835 -783 -739 -749
rect 739 -783 835 -749
<< nsubdiffcont >>
rect -739 749 739 783
rect -835 -687 -801 687
rect 801 -687 835 687
rect -739 -783 739 -749
<< poly >>
rect -675 681 -605 697
rect -675 647 -659 681
rect -621 647 -605 681
rect -675 600 -605 647
rect -547 681 -477 697
rect -547 647 -531 681
rect -493 647 -477 681
rect -547 600 -477 647
rect -419 681 -349 697
rect -419 647 -403 681
rect -365 647 -349 681
rect -419 600 -349 647
rect -291 681 -221 697
rect -291 647 -275 681
rect -237 647 -221 681
rect -291 600 -221 647
rect -163 681 -93 697
rect -163 647 -147 681
rect -109 647 -93 681
rect -163 600 -93 647
rect -35 681 35 697
rect -35 647 -19 681
rect 19 647 35 681
rect -35 600 35 647
rect 93 681 163 697
rect 93 647 109 681
rect 147 647 163 681
rect 93 600 163 647
rect 221 681 291 697
rect 221 647 237 681
rect 275 647 291 681
rect 221 600 291 647
rect 349 681 419 697
rect 349 647 365 681
rect 403 647 419 681
rect 349 600 419 647
rect 477 681 547 697
rect 477 647 493 681
rect 531 647 547 681
rect 477 600 547 647
rect 605 681 675 697
rect 605 647 621 681
rect 659 647 675 681
rect 605 600 675 647
rect -675 -647 -605 -600
rect -675 -681 -659 -647
rect -621 -681 -605 -647
rect -675 -697 -605 -681
rect -547 -647 -477 -600
rect -547 -681 -531 -647
rect -493 -681 -477 -647
rect -547 -697 -477 -681
rect -419 -647 -349 -600
rect -419 -681 -403 -647
rect -365 -681 -349 -647
rect -419 -697 -349 -681
rect -291 -647 -221 -600
rect -291 -681 -275 -647
rect -237 -681 -221 -647
rect -291 -697 -221 -681
rect -163 -647 -93 -600
rect -163 -681 -147 -647
rect -109 -681 -93 -647
rect -163 -697 -93 -681
rect -35 -647 35 -600
rect -35 -681 -19 -647
rect 19 -681 35 -647
rect -35 -697 35 -681
rect 93 -647 163 -600
rect 93 -681 109 -647
rect 147 -681 163 -647
rect 93 -697 163 -681
rect 221 -647 291 -600
rect 221 -681 237 -647
rect 275 -681 291 -647
rect 221 -697 291 -681
rect 349 -647 419 -600
rect 349 -681 365 -647
rect 403 -681 419 -647
rect 349 -697 419 -681
rect 477 -647 547 -600
rect 477 -681 493 -647
rect 531 -681 547 -647
rect 477 -697 547 -681
rect 605 -647 675 -600
rect 605 -681 621 -647
rect 659 -681 675 -647
rect 605 -697 675 -681
<< polycont >>
rect -659 647 -621 681
rect -531 647 -493 681
rect -403 647 -365 681
rect -275 647 -237 681
rect -147 647 -109 681
rect -19 647 19 681
rect 109 647 147 681
rect 237 647 275 681
rect 365 647 403 681
rect 493 647 531 681
rect 621 647 659 681
rect -659 -681 -621 -647
rect -531 -681 -493 -647
rect -403 -681 -365 -647
rect -275 -681 -237 -647
rect -147 -681 -109 -647
rect -19 -681 19 -647
rect 109 -681 147 -647
rect 237 -681 275 -647
rect 365 -681 403 -647
rect 493 -681 531 -647
rect 621 -681 659 -647
<< locali >>
rect -835 749 -739 783
rect 739 749 835 783
rect -835 687 -801 749
rect 801 687 835 749
rect -675 647 -659 681
rect -621 647 -605 681
rect -547 647 -531 681
rect -493 647 -477 681
rect -419 647 -403 681
rect -365 647 -349 681
rect -291 647 -275 681
rect -237 647 -221 681
rect -163 647 -147 681
rect -109 647 -93 681
rect -35 647 -19 681
rect 19 647 35 681
rect 93 647 109 681
rect 147 647 163 681
rect 221 647 237 681
rect 275 647 291 681
rect 349 647 365 681
rect 403 647 419 681
rect 477 647 493 681
rect 531 647 547 681
rect 605 647 621 681
rect 659 647 675 681
rect -721 588 -687 604
rect -721 -604 -687 -588
rect -593 588 -559 604
rect -593 -604 -559 -588
rect -465 588 -431 604
rect -465 -604 -431 -588
rect -337 588 -303 604
rect -337 -604 -303 -588
rect -209 588 -175 604
rect -209 -604 -175 -588
rect -81 588 -47 604
rect -81 -604 -47 -588
rect 47 588 81 604
rect 47 -604 81 -588
rect 175 588 209 604
rect 175 -604 209 -588
rect 303 588 337 604
rect 303 -604 337 -588
rect 431 588 465 604
rect 431 -604 465 -588
rect 559 588 593 604
rect 559 -604 593 -588
rect 687 588 721 604
rect 687 -604 721 -588
rect -675 -681 -659 -647
rect -621 -681 -605 -647
rect -547 -681 -531 -647
rect -493 -681 -477 -647
rect -419 -681 -403 -647
rect -365 -681 -349 -647
rect -291 -681 -275 -647
rect -237 -681 -221 -647
rect -163 -681 -147 -647
rect -109 -681 -93 -647
rect -35 -681 -19 -647
rect 19 -681 35 -647
rect 93 -681 109 -647
rect 147 -681 163 -647
rect 221 -681 237 -647
rect 275 -681 291 -647
rect 349 -681 365 -647
rect 403 -681 419 -647
rect 477 -681 493 -647
rect 531 -681 547 -647
rect 605 -681 621 -647
rect 659 -681 675 -647
rect -835 -749 -801 -687
rect 801 -749 835 -687
rect -835 -783 -739 -749
rect 739 -783 835 -749
<< viali >>
rect -659 647 -621 681
rect -531 647 -493 681
rect -403 647 -365 681
rect -275 647 -237 681
rect -147 647 -109 681
rect -19 647 19 681
rect 109 647 147 681
rect 237 647 275 681
rect 365 647 403 681
rect 493 647 531 681
rect 621 647 659 681
rect -721 -588 -687 588
rect -593 -588 -559 588
rect -465 -588 -431 588
rect -337 -588 -303 588
rect -209 -588 -175 588
rect -81 -588 -47 588
rect 47 -588 81 588
rect 175 -588 209 588
rect 303 -588 337 588
rect 431 -588 465 588
rect 559 -588 593 588
rect 687 -588 721 588
rect -659 -681 -621 -647
rect -531 -681 -493 -647
rect -403 -681 -365 -647
rect -275 -681 -237 -647
rect -147 -681 -109 -647
rect -19 -681 19 -647
rect 109 -681 147 -647
rect 237 -681 275 -647
rect 365 -681 403 -647
rect 493 -681 531 -647
rect 621 -681 659 -647
<< metal1 >>
rect -671 681 -609 687
rect -671 647 -659 681
rect -621 647 -609 681
rect -671 641 -609 647
rect -543 681 -481 687
rect -543 647 -531 681
rect -493 647 -481 681
rect -543 641 -481 647
rect -415 681 -353 687
rect -415 647 -403 681
rect -365 647 -353 681
rect -415 641 -353 647
rect -287 681 -225 687
rect -287 647 -275 681
rect -237 647 -225 681
rect -287 641 -225 647
rect -159 681 -97 687
rect -159 647 -147 681
rect -109 647 -97 681
rect -159 641 -97 647
rect -31 681 31 687
rect -31 647 -19 681
rect 19 647 31 681
rect -31 641 31 647
rect 97 681 159 687
rect 97 647 109 681
rect 147 647 159 681
rect 97 641 159 647
rect 225 681 287 687
rect 225 647 237 681
rect 275 647 287 681
rect 225 641 287 647
rect 353 681 415 687
rect 353 647 365 681
rect 403 647 415 681
rect 353 641 415 647
rect 481 681 543 687
rect 481 647 493 681
rect 531 647 543 681
rect 481 641 543 647
rect 609 681 671 687
rect 609 647 621 681
rect 659 647 671 681
rect 609 641 671 647
rect -727 588 -681 600
rect -727 -588 -721 588
rect -687 -588 -681 588
rect -727 -600 -681 -588
rect -599 588 -553 600
rect -599 -588 -593 588
rect -559 -588 -553 588
rect -599 -600 -553 -588
rect -471 588 -425 600
rect -471 -588 -465 588
rect -431 -588 -425 588
rect -471 -600 -425 -588
rect -343 588 -297 600
rect -343 -588 -337 588
rect -303 -588 -297 588
rect -343 -600 -297 -588
rect -215 588 -169 600
rect -215 -588 -209 588
rect -175 -588 -169 588
rect -215 -600 -169 -588
rect -87 588 -41 600
rect -87 -588 -81 588
rect -47 -588 -41 588
rect -87 -600 -41 -588
rect 41 588 87 600
rect 41 -588 47 588
rect 81 -588 87 588
rect 41 -600 87 -588
rect 169 588 215 600
rect 169 -588 175 588
rect 209 -588 215 588
rect 169 -600 215 -588
rect 297 588 343 600
rect 297 -588 303 588
rect 337 -588 343 588
rect 297 -600 343 -588
rect 425 588 471 600
rect 425 -588 431 588
rect 465 -588 471 588
rect 425 -600 471 -588
rect 553 588 599 600
rect 553 -588 559 588
rect 593 -588 599 588
rect 553 -600 599 -588
rect 681 588 727 600
rect 681 -588 687 588
rect 721 -588 727 588
rect 681 -600 727 -588
rect -671 -647 -609 -641
rect -671 -681 -659 -647
rect -621 -681 -609 -647
rect -671 -687 -609 -681
rect -543 -647 -481 -641
rect -543 -681 -531 -647
rect -493 -681 -481 -647
rect -543 -687 -481 -681
rect -415 -647 -353 -641
rect -415 -681 -403 -647
rect -365 -681 -353 -647
rect -415 -687 -353 -681
rect -287 -647 -225 -641
rect -287 -681 -275 -647
rect -237 -681 -225 -647
rect -287 -687 -225 -681
rect -159 -647 -97 -641
rect -159 -681 -147 -647
rect -109 -681 -97 -647
rect -159 -687 -97 -681
rect -31 -647 31 -641
rect -31 -681 -19 -647
rect 19 -681 31 -647
rect -31 -687 31 -681
rect 97 -647 159 -641
rect 97 -681 109 -647
rect 147 -681 159 -647
rect 97 -687 159 -681
rect 225 -647 287 -641
rect 225 -681 237 -647
rect 275 -681 287 -647
rect 225 -687 287 -681
rect 353 -647 415 -641
rect 353 -681 365 -647
rect 403 -681 415 -647
rect 353 -687 415 -681
rect 481 -647 543 -641
rect 481 -681 493 -647
rect 531 -681 543 -647
rect 481 -687 543 -681
rect 609 -647 671 -641
rect 609 -681 621 -647
rect 659 -681 671 -647
rect 609 -687 671 -681
<< properties >>
string FIXED_BBOX -818 -766 818 766
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 6 l 0.35 m 1 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
