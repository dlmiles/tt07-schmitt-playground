magic
tech sky130A
magscale 1 2
timestamp 1717304205
<< nwell >>
rect 21000 41922 21130 42171
<< locali >>
rect 200 40040 31808 40094
rect 200 39976 8148 40040
rect 10502 39976 31808 40040
rect 200 39894 31808 39976
rect 200 39630 628 39894
rect 18714 39758 31808 39894
rect 18714 39630 31518 39758
rect 200 39553 31518 39630
rect 200 39489 239 39553
rect 200 39488 31518 39489
rect 31772 39488 31808 39758
rect 200 39430 31808 39488
<< viali >>
rect 857 44471 891 44505
rect 1593 44471 1627 44505
rect 2329 44471 2363 44505
rect 3249 44471 3283 44505
rect 3801 44471 3835 44505
rect 4537 44471 4571 44505
rect 5273 44471 5307 44505
rect 6009 44471 6043 44505
rect 14105 44471 14139 44505
rect 15577 44471 15611 44505
rect 18061 44471 18095 44505
rect 19073 44471 19107 44505
rect 23397 44471 23431 44505
rect 27353 44471 27387 44505
rect 28457 44471 28491 44505
rect 11621 44403 11655 44437
rect 12909 44403 12943 44437
rect 17049 44403 17083 44437
rect 24961 44403 24995 44437
rect 29377 44403 29411 44437
rect 30665 44403 30699 44437
rect 11897 44356 11931 44390
rect 12357 44356 12391 44390
rect 13185 44335 13219 44369
rect 13691 44351 13725 44385
rect 13829 44351 13863 44385
rect 14289 44335 14323 44369
rect 15485 44359 15519 44393
rect 15761 44369 15795 44403
rect 16497 44356 16531 44390
rect 16865 44356 16899 44390
rect 18889 44369 18923 44403
rect 17417 44335 17451 44369
rect 19165 44343 19199 44377
rect 19257 44343 19291 44377
rect 21925 44335 21959 44369
rect 22017 44343 22051 44377
rect 22753 44335 22787 44369
rect 23121 44335 23155 44369
rect 23213 44335 23247 44369
rect 24777 44335 24811 44369
rect 25237 44335 25271 44369
rect 25513 44335 25547 44369
rect 26801 44335 26835 44369
rect 27261 44335 27295 44369
rect 27721 44335 27755 44369
rect 28273 44335 28307 44369
rect 28641 44335 28675 44369
rect 30205 44335 30239 44369
rect 31217 44335 31251 44369
rect 12700 44267 12734 44301
rect 12817 44267 12851 44301
rect 24593 44267 24627 44301
rect 25329 44267 25363 44301
rect 27445 44267 27479 44301
rect 29101 44267 29135 44301
rect 29285 44267 29319 44301
rect 29929 44267 29963 44301
rect 30113 44267 30147 44301
rect 12541 44199 12575 44233
rect 13829 44199 13863 44233
rect 15945 44199 15979 44233
rect 18705 44199 18739 44233
rect 19349 44199 19383 44233
rect 21281 44199 21315 44233
rect 22109 44199 22143 44233
rect 25053 44199 25087 44233
rect 26617 44199 26651 44233
rect 26893 44199 26927 44233
rect 29745 44199 29779 44233
rect 30573 44199 30607 44233
rect 15301 43927 15335 43961
rect 17233 43927 17267 43961
rect 21465 43927 21499 43961
rect 23673 43927 23707 43961
rect 30389 43927 30423 43961
rect 30573 43927 30607 43961
rect 21557 43859 21591 43893
rect 10977 43791 11011 43825
rect 11713 43791 11747 43825
rect 13553 43791 13587 43825
rect 15117 43791 15151 43825
rect 15853 43791 15887 43825
rect 17417 43791 17451 43825
rect 18705 43791 18739 43825
rect 22937 43791 22971 43825
rect 28181 43791 28215 43825
rect 31125 43791 31159 43825
rect 10885 43735 10919 43769
rect 11529 43723 11563 43757
rect 11980 43723 12014 43757
rect 13921 43723 13955 43757
rect 14381 43738 14415 43772
rect 14841 43738 14875 43772
rect 15017 43751 15051 43785
rect 15485 43723 15519 43757
rect 15761 43723 15795 43757
rect 16120 43723 16154 43757
rect 17601 43738 17635 43772
rect 17877 43738 17911 43772
rect 19349 43723 19383 43757
rect 19625 43723 19659 43757
rect 19901 43723 19935 43757
rect 20085 43723 20119 43757
rect 20352 43723 20386 43757
rect 22670 43723 22704 43757
rect 23397 43723 23431 43757
rect 23489 43723 23523 43757
rect 24041 43735 24075 43769
rect 24317 43723 24351 43757
rect 24562 43723 24596 43757
rect 26617 43723 26651 43757
rect 26884 43723 26918 43757
rect 29009 43723 29043 43757
rect 29276 43723 29310 43757
rect 11253 43655 11287 43689
rect 13093 43655 13127 43689
rect 14749 43655 14783 43689
rect 15669 43655 15703 43689
rect 19441 43655 19475 43689
rect 19809 43655 19843 43689
rect 23029 43655 23063 43689
rect 23949 43655 23983 43689
rect 25697 43655 25731 43689
rect 27997 43655 28031 43689
rect 28365 43655 28399 43689
rect 28457 43655 28491 43689
rect 28825 43655 28859 43689
rect 14197 43383 14231 43417
rect 14473 43383 14507 43417
rect 22937 43383 22971 43417
rect 25973 43383 26007 43417
rect 26893 43383 26927 43417
rect 28917 43383 28951 43417
rect 29193 43383 29227 43417
rect 30941 43383 30975 43417
rect 19625 43349 19659 43383
rect 13185 43315 13219 43349
rect 16396 43315 16430 43349
rect 18806 43315 18840 43349
rect 23826 43315 23860 43349
rect 25145 43315 25179 43349
rect 25513 43315 25547 43349
rect 28580 43315 28614 43349
rect 29736 43315 29770 43349
rect 13093 43247 13127 43281
rect 14356 43247 14390 43281
rect 14841 43247 14875 43281
rect 15025 43267 15059 43301
rect 15753 43255 15787 43289
rect 15853 43247 15887 43281
rect 16129 43247 16163 43281
rect 19073 43247 19107 43281
rect 19349 43247 19383 43281
rect 21465 43247 21499 43281
rect 23581 43247 23615 43281
rect 25237 43255 25271 43289
rect 26617 43247 26651 43281
rect 27077 43247 27111 43281
rect 28825 43247 28859 43281
rect 29101 43247 29135 43281
rect 29377 43247 29411 43281
rect 29469 43247 29503 43281
rect 31125 43247 31159 43281
rect 11345 43179 11379 43213
rect 13461 43179 13495 43213
rect 14565 43179 14599 43213
rect 17693 43179 17727 43213
rect 24961 43179 24995 43213
rect 26065 43179 26099 43213
rect 26249 43179 26283 43213
rect 27445 43179 27479 43213
rect 25513 43145 25547 43179
rect 15209 43111 15243 43145
rect 17509 43111 17543 43145
rect 21097 43111 21131 43145
rect 26433 43111 26467 43145
rect 30849 43111 30883 43145
rect 11161 42839 11195 42873
rect 11713 42839 11747 42873
rect 16865 42839 16899 42873
rect 23397 42839 23431 42873
rect 28641 42839 28675 42873
rect 29193 42839 29227 42873
rect 29285 42839 29319 42873
rect 30481 42839 30515 42873
rect 12725 42771 12759 42805
rect 24041 42771 24075 42805
rect 15209 42737 15243 42771
rect 11989 42703 12023 42737
rect 12265 42703 12299 42737
rect 14749 42703 14783 42737
rect 21005 42703 21039 42737
rect 21281 42703 21315 42737
rect 21833 42703 21867 42737
rect 22569 42703 22603 42737
rect 23121 42703 23155 42737
rect 24409 42703 24443 42737
rect 26433 42703 26467 42737
rect 27997 42703 28031 42737
rect 11253 42635 11287 42669
rect 11805 42635 11839 42669
rect 13001 42635 13035 42669
rect 13369 42635 13403 42669
rect 13691 42650 13725 42684
rect 14289 42650 14323 42684
rect 15301 42635 15335 42669
rect 15577 42635 15611 42669
rect 15853 42650 15887 42684
rect 16313 42650 16347 42684
rect 18153 42635 18187 42669
rect 18429 42635 18463 42669
rect 23213 42635 23247 42669
rect 23673 42635 23707 42669
rect 24317 42635 24351 42669
rect 24676 42635 24710 42669
rect 26617 42635 26651 42669
rect 26801 42635 26835 42669
rect 29009 42635 29043 42669
rect 29469 42635 29503 42669
rect 30665 42635 30699 42669
rect 12725 42601 12759 42635
rect 12173 42567 12207 42601
rect 14197 42567 14231 42601
rect 14933 42567 14967 42601
rect 18245 42567 18279 42601
rect 20453 42567 20487 42601
rect 20821 42567 20855 42601
rect 20913 42567 20947 42601
rect 22017 42567 22051 42601
rect 22753 42567 22787 42601
rect 23489 42567 23523 42601
rect 23857 42567 23891 42601
rect 25789 42567 25823 42601
rect 25881 42567 25915 42601
rect 12081 42295 12115 42329
rect 12357 42295 12391 42329
rect 13185 42295 13219 42329
rect 22109 42295 22143 42329
rect 22753 42295 22787 42329
rect 23397 42295 23431 42329
rect 2982 42227 3016 42261
rect 11805 42227 11839 42261
rect 12265 42227 12299 42261
rect 12817 42227 12851 42261
rect 20269 42227 20303 42261
rect 22293 42227 22327 42261
rect 14565 42193 14599 42227
rect 3249 42159 3283 42193
rect 3433 42159 3467 42193
rect 13001 42159 13035 42193
rect 13480 42159 13514 42193
rect 13578 42159 13612 42193
rect 14105 42159 14139 42193
rect 14381 42159 14415 42193
rect 15209 42180 15243 42214
rect 15669 42180 15703 42214
rect 16313 42159 16347 42193
rect 17048 42175 17082 42209
rect 17233 42159 17267 42193
rect 17325 42183 17359 42217
rect 20085 42193 20119 42227
rect 21465 42193 21499 42227
rect 21649 42193 21683 42227
rect 21751 42193 21785 42227
rect 19625 42159 19659 42193
rect 20453 42159 20487 42193
rect 20637 42159 20671 42193
rect 20729 42159 20763 42193
rect 22385 42175 22419 42209
rect 22569 42175 22603 42209
rect 24757 42193 24791 42227
rect 23121 42159 23155 42193
rect 23213 42159 23247 42193
rect 24501 42159 24535 42193
rect 26985 42159 27019 42193
rect 11437 42091 11471 42125
rect 14749 42091 14783 42125
rect 15669 42091 15703 42125
rect 16497 42091 16531 42125
rect 16865 42091 16899 42125
rect 19441 42091 19475 42125
rect 19809 42091 19843 42125
rect 21281 42091 21315 42125
rect 25881 42091 25915 42125
rect 12817 42057 12851 42091
rect 1869 42023 1903 42057
rect 4077 42023 4111 42057
rect 11989 42023 12023 42057
rect 16129 42023 16163 42057
rect 19901 42023 19935 42057
rect 20913 42023 20947 42057
rect 21925 42023 21959 42057
rect 22569 42023 22603 42057
rect 26433 42023 26467 42057
rect 11805 41973 11839 42007
rect 14289 41973 14323 42007
rect 22143 41973 22177 42007
rect 14197 41751 14231 41785
rect 21603 41751 21637 41785
rect 25697 41761 25731 41795
rect 25881 41751 25915 41785
rect 6653 41683 6687 41717
rect 22385 41683 22419 41717
rect 16405 41649 16439 41683
rect 2421 41615 2455 41649
rect 6009 41615 6043 41649
rect 15393 41615 15427 41649
rect 16313 41615 16347 41649
rect 16865 41615 16899 41649
rect 16957 41615 16991 41649
rect 17969 41615 18003 41649
rect 19257 41615 19291 41649
rect 19717 41615 19751 41649
rect 22201 41615 22235 41649
rect 2329 41547 2363 41581
rect 3893 41547 3927 41581
rect 4160 41547 4194 41581
rect 11713 41547 11747 41581
rect 12035 41562 12069 41596
rect 12449 41562 12483 41596
rect 12817 41562 12851 41596
rect 13001 41562 13035 41596
rect 13737 41575 13771 41609
rect 14105 41562 14139 41596
rect 15117 41564 15151 41598
rect 15563 41559 15597 41593
rect 17141 41559 17175 41593
rect 18139 41559 18173 41593
rect 19441 41581 19475 41615
rect 22014 41581 22048 41615
rect 22477 41562 22511 41596
rect 22661 41562 22695 41596
rect 25421 41575 25455 41609
rect 3065 41479 3099 41513
rect 5273 41479 5307 41513
rect 13185 41479 13219 41513
rect 13645 41479 13679 41513
rect 15761 41479 15795 41513
rect 16681 41479 16715 41513
rect 17325 41479 17359 41513
rect 18337 41479 18371 41513
rect 19625 41479 19659 41513
rect 19993 41479 20027 41513
rect 21833 41479 21867 41513
rect 2145 41207 2179 41241
rect 2513 41207 2547 41241
rect 4353 41207 4387 41241
rect 6561 41207 6595 41241
rect 8033 41207 8067 41241
rect 11805 41207 11839 41241
rect 15669 41207 15703 41241
rect 17969 41207 18003 41241
rect 20453 41207 20487 41241
rect 22201 41207 22235 41241
rect 3626 41139 3660 41173
rect 14289 41139 14323 41173
rect 17693 41139 17727 41173
rect 19257 41139 19291 41173
rect 20729 41139 20763 41173
rect 21833 41139 21867 41173
rect 30205 41139 30239 41173
rect 2329 41071 2363 41105
rect 3893 41071 3927 41105
rect 4537 41071 4571 41105
rect 6745 41071 6779 41105
rect 8217 41071 8251 41105
rect 11989 41092 12023 41126
rect 12173 41092 12207 41126
rect 12541 41071 12575 41105
rect 12650 41071 12684 41105
rect 12817 41092 12851 41126
rect 13645 41091 13679 41125
rect 14104 41105 14138 41139
rect 14381 41071 14415 41105
rect 14565 41092 14599 41126
rect 15117 41092 15151 41126
rect 15347 41092 15381 41126
rect 15945 41092 15979 41126
rect 16405 41092 16439 41126
rect 16589 41092 16623 41126
rect 16957 41092 16991 41126
rect 17371 41092 17405 41126
rect 17785 41071 17819 41105
rect 20269 41071 20303 41105
rect 22017 41071 22051 41105
rect 23481 41095 23515 41129
rect 23581 41071 23615 41105
rect 30492 41088 30526 41122
rect 13829 41003 13863 41037
rect 16129 41003 16163 41037
rect 21005 41003 21039 41037
rect 19533 40935 19567 40969
rect 21741 40935 21775 40969
rect 13093 40527 13127 40561
rect 12889 40471 12923 40505
rect 15025 40459 15059 40493
rect 15209 40474 15243 40508
rect 15669 40474 15703 40508
rect 16129 40459 16163 40493
rect 12725 40391 12759 40425
rect 16313 40391 16347 40425
rect 8148 39976 10502 40040
rect 31518 39553 31772 39758
rect 239 39489 31772 39553
rect 31518 39488 31772 39489
<< metal1 >>
rect 15746 44734 15752 44786
rect 15804 44774 15810 44786
rect 23290 44774 23296 44786
rect 15804 44746 23296 44774
rect 15804 44734 15810 44746
rect 23290 44734 23296 44746
rect 23348 44734 23354 44786
rect 23474 44734 23480 44786
rect 23532 44774 23538 44786
rect 30374 44774 30380 44786
rect 23532 44746 30380 44774
rect 23532 44734 23538 44746
rect 30374 44734 30380 44746
rect 30432 44734 30438 44786
rect 552 44634 31808 44656
rect 552 44582 8172 44634
rect 8224 44582 8236 44634
rect 8288 44582 8300 44634
rect 8352 44582 8364 44634
rect 8416 44582 8428 44634
rect 8480 44582 15946 44634
rect 15998 44582 16010 44634
rect 16062 44582 16074 44634
rect 16126 44582 16138 44634
rect 16190 44582 16202 44634
rect 16254 44582 23720 44634
rect 23772 44582 23784 44634
rect 23836 44582 23848 44634
rect 23900 44582 23912 44634
rect 23964 44582 23976 44634
rect 24028 44582 31494 44634
rect 31546 44582 31558 44634
rect 31610 44582 31622 44634
rect 31674 44582 31686 44634
rect 31738 44582 31750 44634
rect 31802 44582 31808 44634
rect 552 44560 31808 44582
rect 842 44462 848 44514
rect 900 44462 906 44514
rect 1578 44462 1584 44514
rect 1636 44462 1642 44514
rect 2314 44462 2320 44514
rect 2372 44462 2378 44514
rect 3234 44462 3240 44514
rect 3292 44462 3298 44514
rect 3786 44462 3792 44514
rect 3844 44462 3850 44514
rect 4522 44462 4528 44514
rect 4580 44462 4586 44514
rect 5258 44462 5264 44514
rect 5316 44462 5322 44514
rect 5994 44462 6000 44514
rect 6052 44462 6058 44514
rect 13906 44502 13912 44514
rect 11900 44474 13912 44502
rect 9674 44394 9680 44446
rect 9732 44434 9738 44446
rect 11609 44437 11667 44443
rect 11609 44434 11621 44437
rect 9732 44406 11621 44434
rect 9732 44394 9738 44406
rect 11609 44403 11621 44406
rect 11655 44403 11667 44437
rect 11609 44397 11667 44403
rect 11900 44396 11928 44474
rect 13906 44462 13912 44474
rect 13964 44502 13970 44514
rect 13964 44474 14044 44502
rect 13964 44462 13970 44474
rect 12897 44437 12955 44443
rect 12897 44403 12909 44437
rect 12943 44434 12955 44437
rect 13354 44434 13360 44446
rect 12943 44406 13360 44434
rect 12943 44403 12955 44406
rect 11885 44390 11943 44396
rect 11885 44356 11897 44390
rect 11931 44356 11943 44390
rect 11885 44350 11943 44356
rect 12345 44390 12403 44396
rect 12345 44356 12357 44390
rect 12391 44387 12403 44390
rect 12618 44387 12624 44399
rect 12391 44359 12624 44387
rect 12391 44356 12403 44359
rect 12345 44350 12403 44356
rect 12618 44347 12624 44359
rect 12676 44347 12682 44399
rect 12897 44397 12955 44403
rect 13354 44394 13360 44406
rect 13412 44394 13418 44446
rect 14016 44434 14044 44474
rect 14090 44462 14096 44514
rect 14148 44462 14154 44514
rect 15565 44505 15623 44511
rect 15565 44471 15577 44505
rect 15611 44502 15623 44505
rect 15654 44502 15660 44514
rect 15611 44474 15660 44502
rect 15611 44471 15623 44474
rect 15565 44465 15623 44471
rect 15654 44462 15660 44474
rect 15712 44462 15718 44514
rect 17862 44502 17868 44514
rect 16592 44474 17868 44502
rect 14366 44434 14372 44446
rect 14016 44406 14372 44434
rect 14366 44394 14372 44406
rect 14424 44394 14430 44446
rect 13679 44385 13737 44391
rect 13173 44369 13231 44375
rect 13173 44335 13185 44369
rect 13219 44366 13231 44369
rect 13538 44366 13544 44378
rect 13219 44338 13544 44366
rect 13219 44335 13231 44338
rect 13173 44329 13231 44335
rect 13538 44326 13544 44338
rect 13596 44326 13602 44378
rect 13679 44351 13691 44385
rect 13725 44351 13737 44385
rect 13679 44345 13737 44351
rect 12688 44301 12746 44307
rect 12688 44267 12700 44301
rect 12734 44298 12746 44301
rect 12805 44301 12863 44307
rect 12734 44267 12756 44298
rect 12688 44261 12756 44267
rect 12805 44267 12817 44301
rect 12851 44298 12863 44301
rect 13262 44298 13268 44310
rect 12851 44270 13268 44298
rect 12851 44267 12863 44270
rect 12805 44261 12863 44267
rect 12526 44190 12532 44242
rect 12584 44190 12590 44242
rect 12728 44230 12756 44261
rect 13262 44258 13268 44270
rect 13320 44258 13326 44310
rect 13354 44258 13360 44310
rect 13412 44298 13418 44310
rect 13694 44298 13722 44345
rect 13814 44342 13820 44394
rect 13872 44342 13878 44394
rect 15473 44393 15531 44399
rect 14274 44326 14280 44378
rect 14332 44326 14338 44378
rect 15473 44359 15485 44393
rect 15519 44390 15531 44393
rect 15562 44390 15568 44402
rect 15519 44362 15568 44390
rect 15519 44359 15531 44362
rect 15473 44353 15531 44359
rect 15562 44350 15568 44362
rect 15620 44350 15626 44402
rect 15746 44360 15752 44412
rect 15804 44360 15810 44412
rect 16298 44347 16304 44399
rect 16356 44387 16362 44399
rect 16485 44390 16543 44396
rect 16485 44387 16497 44390
rect 16356 44359 16497 44387
rect 16356 44347 16362 44359
rect 16485 44356 16497 44359
rect 16531 44387 16543 44390
rect 16592 44387 16620 44474
rect 17862 44462 17868 44474
rect 17920 44462 17926 44514
rect 18049 44505 18107 44511
rect 18049 44471 18061 44505
rect 18095 44502 18107 44505
rect 19061 44505 19119 44511
rect 19061 44502 19073 44505
rect 18095 44474 19073 44502
rect 18095 44471 18107 44474
rect 18049 44465 18107 44471
rect 19061 44471 19073 44474
rect 19107 44471 19119 44505
rect 19061 44465 19119 44471
rect 19150 44462 19156 44514
rect 19208 44502 19214 44514
rect 19208 44474 19564 44502
rect 19208 44462 19214 44474
rect 16531 44359 16620 44387
rect 16531 44356 16543 44359
rect 16485 44350 16543 44356
rect 16850 44347 16856 44399
rect 16908 44347 16914 44399
rect 17034 44394 17040 44446
rect 17092 44394 17098 44446
rect 19536 44434 19564 44474
rect 19610 44462 19616 44514
rect 19668 44502 19674 44514
rect 23385 44505 23443 44511
rect 23385 44502 23397 44505
rect 19668 44474 23397 44502
rect 19668 44462 19674 44474
rect 23385 44471 23397 44474
rect 23431 44471 23443 44505
rect 27341 44505 27399 44511
rect 23385 44465 23443 44471
rect 24872 44474 27292 44502
rect 21818 44434 21824 44446
rect 18877 44403 18935 44409
rect 19536 44406 21824 44434
rect 17218 44326 17224 44378
rect 17276 44366 17282 44378
rect 17405 44369 17463 44375
rect 17405 44366 17417 44369
rect 17276 44338 17417 44366
rect 17276 44326 17282 44338
rect 17405 44335 17417 44338
rect 17451 44335 17463 44369
rect 18877 44369 18889 44403
rect 18923 44369 18935 44403
rect 21818 44394 21824 44406
rect 21876 44394 21882 44446
rect 24872 44434 24900 44474
rect 23124 44406 24900 44434
rect 24949 44437 25007 44443
rect 18877 44366 18935 44369
rect 18966 44366 18972 44378
rect 18877 44363 18972 44366
rect 18892 44338 18972 44363
rect 17405 44329 17463 44335
rect 18966 44326 18972 44338
rect 19024 44326 19030 44378
rect 19058 44334 19064 44386
rect 19116 44374 19122 44386
rect 19153 44377 19211 44383
rect 19153 44374 19165 44377
rect 19116 44346 19165 44374
rect 19116 44334 19122 44346
rect 19153 44343 19165 44346
rect 19199 44343 19211 44377
rect 19153 44337 19211 44343
rect 19242 44334 19248 44386
rect 19300 44334 19306 44386
rect 21910 44326 21916 44378
rect 21968 44326 21974 44378
rect 22005 44377 22063 44383
rect 22005 44343 22017 44377
rect 22051 44343 22063 44377
rect 22005 44337 22063 44343
rect 14918 44298 14924 44310
rect 13412 44270 14924 44298
rect 13412 44258 13418 44270
rect 14918 44258 14924 44270
rect 14976 44258 14982 44310
rect 15470 44258 15476 44310
rect 15528 44298 15534 44310
rect 21726 44298 21732 44310
rect 15528 44270 21732 44298
rect 15528 44258 15534 44270
rect 21726 44258 21732 44270
rect 21784 44258 21790 44310
rect 22020 44242 22048 44337
rect 22094 44326 22100 44378
rect 22152 44366 22158 44378
rect 22741 44369 22799 44375
rect 22741 44366 22753 44369
rect 22152 44338 22753 44366
rect 22152 44326 22158 44338
rect 22741 44335 22753 44338
rect 22787 44366 22799 44369
rect 23014 44366 23020 44378
rect 22787 44338 23020 44366
rect 22787 44335 22799 44338
rect 22741 44329 22799 44335
rect 23014 44326 23020 44338
rect 23072 44326 23078 44378
rect 23124 44375 23152 44406
rect 24949 44403 24961 44437
rect 24995 44434 25007 44437
rect 26510 44434 26516 44446
rect 24995 44406 26516 44434
rect 24995 44403 25007 44406
rect 24949 44397 25007 44403
rect 26510 44394 26516 44406
rect 26568 44394 26574 44446
rect 27264 44434 27292 44474
rect 27341 44471 27353 44505
rect 27387 44502 27399 44505
rect 28445 44505 28503 44511
rect 28445 44502 28457 44505
rect 27387 44474 28457 44502
rect 27387 44471 27399 44474
rect 27341 44465 27399 44471
rect 28445 44471 28457 44474
rect 28491 44471 28503 44505
rect 31110 44502 31116 44514
rect 28445 44465 28503 44471
rect 29288 44474 31116 44502
rect 29288 44434 29316 44474
rect 31110 44462 31116 44474
rect 31168 44462 31174 44514
rect 27264 44406 29316 44434
rect 29365 44437 29423 44443
rect 29365 44403 29377 44437
rect 29411 44434 29423 44437
rect 30653 44437 30711 44443
rect 30653 44434 30665 44437
rect 29411 44406 30665 44434
rect 29411 44403 29423 44406
rect 29365 44397 29423 44403
rect 30653 44403 30665 44406
rect 30699 44403 30711 44437
rect 30653 44397 30711 44403
rect 23109 44369 23167 44375
rect 23109 44335 23121 44369
rect 23155 44335 23167 44369
rect 23109 44329 23167 44335
rect 23198 44326 23204 44378
rect 23256 44326 23262 44378
rect 24765 44369 24823 44375
rect 24765 44335 24777 44369
rect 24811 44335 24823 44369
rect 24765 44329 24823 44335
rect 24118 44258 24124 44310
rect 24176 44298 24182 44310
rect 24581 44301 24639 44307
rect 24581 44298 24593 44301
rect 24176 44270 24593 44298
rect 24176 44258 24182 44270
rect 24581 44267 24593 44270
rect 24627 44267 24639 44301
rect 24780 44298 24808 44329
rect 25222 44326 25228 44378
rect 25280 44326 25286 44378
rect 25498 44326 25504 44378
rect 25556 44326 25562 44378
rect 26786 44326 26792 44378
rect 26844 44326 26850 44378
rect 27249 44369 27307 44375
rect 27249 44335 27261 44369
rect 27295 44366 27307 44369
rect 27709 44369 27767 44375
rect 27709 44366 27721 44369
rect 27295 44338 27721 44366
rect 27295 44335 27307 44338
rect 27249 44329 27307 44335
rect 27709 44335 27721 44338
rect 27755 44335 27767 44369
rect 27709 44329 27767 44335
rect 27982 44326 27988 44378
rect 28040 44366 28046 44378
rect 28261 44369 28319 44375
rect 28261 44366 28273 44369
rect 28040 44338 28273 44366
rect 28040 44326 28046 44338
rect 28261 44335 28273 44338
rect 28307 44335 28319 44369
rect 28261 44329 28319 44335
rect 28626 44326 28632 44378
rect 28684 44326 28690 44378
rect 30193 44369 30251 44375
rect 29104 44338 29960 44366
rect 25317 44301 25375 44307
rect 25317 44298 25329 44301
rect 24780 44270 25329 44298
rect 24581 44261 24639 44267
rect 25317 44267 25329 44270
rect 25363 44267 25375 44301
rect 25317 44261 25375 44267
rect 13170 44230 13176 44242
rect 12728 44202 13176 44230
rect 13170 44190 13176 44202
rect 13228 44190 13234 44242
rect 13814 44190 13820 44242
rect 13872 44190 13878 44242
rect 15933 44233 15991 44239
rect 15933 44199 15945 44233
rect 15979 44230 15991 44233
rect 16390 44230 16396 44242
rect 15979 44202 16396 44230
rect 15979 44199 15991 44202
rect 15933 44193 15991 44199
rect 16390 44190 16396 44202
rect 16448 44190 16454 44242
rect 16574 44190 16580 44242
rect 16632 44230 16638 44242
rect 18693 44233 18751 44239
rect 18693 44230 18705 44233
rect 16632 44202 18705 44230
rect 16632 44190 16638 44202
rect 18693 44199 18705 44202
rect 18739 44199 18751 44233
rect 18693 44193 18751 44199
rect 19334 44190 19340 44242
rect 19392 44190 19398 44242
rect 21269 44233 21327 44239
rect 21269 44199 21281 44233
rect 21315 44230 21327 44233
rect 21634 44230 21640 44242
rect 21315 44202 21640 44230
rect 21315 44199 21327 44202
rect 21269 44193 21327 44199
rect 21634 44190 21640 44202
rect 21692 44190 21698 44242
rect 22002 44190 22008 44242
rect 22060 44190 22066 44242
rect 22094 44190 22100 44242
rect 22152 44190 22158 44242
rect 24596 44230 24624 44261
rect 26234 44258 26240 44310
rect 26292 44298 26298 44310
rect 27433 44301 27491 44307
rect 27433 44298 27445 44301
rect 26292 44270 27445 44298
rect 26292 44258 26298 44270
rect 27433 44267 27445 44270
rect 27479 44298 27491 44301
rect 27522 44298 27528 44310
rect 27479 44270 27528 44298
rect 27479 44267 27491 44270
rect 27433 44261 27491 44267
rect 27522 44258 27528 44270
rect 27580 44298 27586 44310
rect 29104 44307 29132 44338
rect 29089 44301 29147 44307
rect 29089 44298 29101 44301
rect 27580 44270 29101 44298
rect 27580 44258 27586 44270
rect 29089 44267 29101 44270
rect 29135 44267 29147 44301
rect 29089 44261 29147 44267
rect 29178 44258 29184 44310
rect 29236 44298 29242 44310
rect 29932 44307 29960 44338
rect 30193 44335 30205 44369
rect 30239 44366 30251 44369
rect 30466 44366 30472 44378
rect 30239 44338 30472 44366
rect 30239 44335 30251 44338
rect 30193 44329 30251 44335
rect 30466 44326 30472 44338
rect 30524 44326 30530 44378
rect 30558 44326 30564 44378
rect 30616 44366 30622 44378
rect 31205 44369 31263 44375
rect 31205 44366 31217 44369
rect 30616 44338 31217 44366
rect 30616 44326 30622 44338
rect 31205 44335 31217 44338
rect 31251 44335 31263 44369
rect 31205 44329 31263 44335
rect 29273 44301 29331 44307
rect 29273 44298 29285 44301
rect 29236 44270 29285 44298
rect 29236 44258 29242 44270
rect 29273 44267 29285 44270
rect 29319 44267 29331 44301
rect 29273 44261 29331 44267
rect 29917 44301 29975 44307
rect 29917 44267 29929 44301
rect 29963 44267 29975 44301
rect 29917 44261 29975 44267
rect 30101 44301 30159 44307
rect 30101 44267 30113 44301
rect 30147 44298 30159 44301
rect 30834 44298 30840 44310
rect 30147 44270 30840 44298
rect 30147 44267 30159 44270
rect 30101 44261 30159 44267
rect 30834 44258 30840 44270
rect 30892 44258 30898 44310
rect 25041 44233 25099 44239
rect 25041 44230 25053 44233
rect 24596 44202 25053 44230
rect 25041 44199 25053 44202
rect 25087 44199 25099 44233
rect 25041 44193 25099 44199
rect 26602 44190 26608 44242
rect 26660 44190 26666 44242
rect 26881 44233 26939 44239
rect 26881 44199 26893 44233
rect 26927 44230 26939 44233
rect 27062 44230 27068 44242
rect 26927 44202 27068 44230
rect 26927 44199 26939 44202
rect 26881 44193 26939 44199
rect 27062 44190 27068 44202
rect 27120 44190 27126 44242
rect 29454 44190 29460 44242
rect 29512 44230 29518 44242
rect 29733 44233 29791 44239
rect 29733 44230 29745 44233
rect 29512 44202 29745 44230
rect 29512 44190 29518 44202
rect 29733 44199 29745 44202
rect 29779 44199 29791 44233
rect 29733 44193 29791 44199
rect 30558 44190 30564 44242
rect 30616 44190 30622 44242
rect 200 44090 31648 44112
rect 200 44038 206 44090
rect 514 44038 4285 44090
rect 4337 44038 4349 44090
rect 4401 44038 4413 44090
rect 4465 44038 4477 44090
rect 4529 44038 4541 44090
rect 4593 44038 12059 44090
rect 12111 44038 12123 44090
rect 12175 44038 12187 44090
rect 12239 44038 12251 44090
rect 12303 44038 12315 44090
rect 12367 44038 19833 44090
rect 19885 44038 19897 44090
rect 19949 44038 19961 44090
rect 20013 44038 20025 44090
rect 20077 44038 20089 44090
rect 20141 44038 27607 44090
rect 27659 44038 27671 44090
rect 27723 44038 27735 44090
rect 27787 44038 27799 44090
rect 27851 44038 27863 44090
rect 27915 44038 31648 44090
rect 200 44016 31648 44038
rect 15289 43961 15347 43967
rect 15289 43958 15301 43961
rect 12912 43930 15301 43958
rect 10965 43825 11023 43831
rect 10965 43791 10977 43825
rect 11011 43822 11023 43825
rect 11701 43825 11759 43831
rect 11701 43822 11713 43825
rect 11011 43794 11713 43822
rect 11011 43791 11023 43794
rect 10965 43785 11023 43791
rect 11701 43791 11713 43794
rect 11747 43791 11759 43825
rect 11701 43785 11759 43791
rect 10873 43769 10931 43775
rect 10873 43735 10885 43769
rect 10919 43754 10931 43769
rect 11330 43754 11336 43766
rect 10919 43735 11336 43754
rect 10873 43729 11336 43735
rect 10888 43726 11336 43729
rect 11330 43714 11336 43726
rect 11388 43714 11394 43766
rect 11514 43714 11520 43766
rect 11572 43714 11578 43766
rect 11968 43757 12026 43763
rect 11968 43723 11980 43757
rect 12014 43754 12026 43757
rect 12912 43754 12940 43930
rect 15289 43927 15301 43930
rect 15335 43927 15347 43961
rect 15289 43921 15347 43927
rect 17218 43918 17224 43970
rect 17276 43918 17282 43970
rect 21453 43961 21511 43967
rect 21453 43927 21465 43961
rect 21499 43958 21511 43961
rect 22002 43958 22008 43970
rect 21499 43930 22008 43958
rect 21499 43927 21511 43930
rect 21453 43921 21511 43927
rect 22002 43918 22008 43930
rect 22060 43918 22066 43970
rect 23658 43918 23664 43970
rect 23716 43918 23722 43970
rect 27522 43918 27528 43970
rect 27580 43958 27586 43970
rect 27580 43930 28028 43958
rect 27580 43918 27586 43930
rect 19058 43890 19064 43902
rect 12014 43726 12940 43754
rect 13004 43862 15048 43890
rect 12014 43723 12026 43726
rect 11968 43717 12026 43723
rect 11238 43646 11244 43698
rect 11296 43646 11302 43698
rect 11348 43686 11376 43714
rect 13004 43686 13032 43862
rect 13541 43825 13599 43831
rect 13541 43791 13553 43825
rect 13587 43822 13599 43825
rect 13998 43822 14004 43834
rect 13587 43794 14004 43822
rect 13587 43791 13599 43794
rect 13541 43785 13599 43791
rect 13998 43782 14004 43794
rect 14056 43782 14062 43834
rect 15020 43791 15048 43862
rect 16863 43862 19064 43890
rect 15105 43825 15163 43831
rect 15105 43791 15117 43825
rect 15151 43822 15163 43825
rect 15841 43825 15899 43831
rect 15841 43822 15853 43825
rect 15151 43794 15853 43822
rect 15151 43791 15163 43794
rect 15005 43785 15063 43791
rect 15105 43785 15163 43791
rect 15841 43791 15853 43794
rect 15887 43791 15899 43825
rect 15841 43785 15899 43791
rect 13909 43757 13967 43763
rect 13909 43723 13921 43757
rect 13955 43754 13967 43757
rect 14182 43754 14188 43766
rect 13955 43726 14188 43754
rect 13955 43723 13967 43726
rect 13909 43717 13967 43723
rect 14182 43714 14188 43726
rect 14240 43714 14246 43766
rect 14366 43729 14372 43781
rect 14424 43729 14430 43781
rect 14829 43772 14887 43778
rect 14829 43738 14841 43772
rect 14875 43738 14887 43772
rect 15005 43751 15017 43785
rect 15051 43754 15063 43785
rect 15378 43754 15384 43766
rect 15051 43751 15384 43754
rect 15005 43745 15384 43751
rect 14829 43732 14887 43738
rect 11348 43658 13032 43686
rect 13081 43689 13139 43695
rect 13081 43655 13093 43689
rect 13127 43686 13139 43689
rect 13170 43686 13176 43698
rect 13127 43658 13176 43686
rect 13127 43655 13139 43658
rect 13081 43649 13139 43655
rect 13170 43646 13176 43658
rect 13228 43646 13234 43698
rect 13998 43646 14004 43698
rect 14056 43686 14062 43698
rect 14458 43686 14464 43698
rect 14056 43658 14464 43686
rect 14056 43646 14062 43658
rect 14458 43646 14464 43658
rect 14516 43646 14522 43698
rect 14734 43646 14740 43698
rect 14792 43646 14798 43698
rect 14844 43686 14872 43732
rect 15020 43726 15384 43745
rect 15378 43714 15384 43726
rect 15436 43714 15442 43766
rect 15470 43714 15476 43766
rect 15528 43714 15534 43766
rect 15562 43714 15568 43766
rect 15620 43754 15626 43766
rect 15749 43757 15807 43763
rect 15749 43754 15761 43757
rect 15620 43726 15761 43754
rect 15620 43714 15626 43726
rect 15749 43723 15761 43726
rect 15795 43723 15807 43757
rect 15749 43717 15807 43723
rect 16108 43757 16166 43763
rect 16108 43723 16120 43757
rect 16154 43754 16166 43757
rect 16574 43754 16580 43766
rect 16154 43726 16580 43754
rect 16154 43723 16166 43726
rect 16108 43717 16166 43723
rect 15194 43686 15200 43698
rect 14844 43658 15200 43686
rect 15194 43646 15200 43658
rect 15252 43646 15258 43698
rect 15286 43646 15292 43698
rect 15344 43686 15350 43698
rect 15657 43689 15715 43695
rect 15657 43686 15669 43689
rect 15344 43658 15669 43686
rect 15344 43646 15350 43658
rect 15657 43655 15669 43658
rect 15703 43655 15715 43689
rect 15764 43686 15792 43717
rect 16574 43714 16580 43726
rect 16632 43714 16638 43766
rect 16863 43686 16891 43862
rect 19058 43850 19064 43862
rect 19116 43890 19122 43902
rect 19886 43890 19892 43902
rect 19116 43862 19892 43890
rect 19116 43850 19122 43862
rect 19886 43850 19892 43862
rect 19944 43850 19950 43902
rect 21545 43893 21603 43899
rect 21545 43859 21557 43893
rect 21591 43890 21603 43893
rect 21910 43890 21916 43902
rect 21591 43862 21916 43890
rect 21591 43859 21603 43862
rect 21545 43853 21603 43859
rect 21910 43850 21916 43862
rect 21968 43850 21974 43902
rect 23198 43850 23204 43902
rect 23256 43890 23262 43902
rect 28000 43890 28028 43930
rect 28074 43918 28080 43970
rect 28132 43958 28138 43970
rect 28902 43958 28908 43970
rect 28132 43930 28908 43958
rect 28132 43918 28138 43930
rect 28902 43918 28908 43930
rect 28960 43918 28966 43970
rect 30374 43918 30380 43970
rect 30432 43918 30438 43970
rect 30466 43918 30472 43970
rect 30524 43958 30530 43970
rect 30561 43961 30619 43967
rect 30561 43958 30573 43961
rect 30524 43930 30573 43958
rect 30524 43918 30530 43930
rect 30561 43927 30573 43930
rect 30607 43927 30619 43961
rect 30561 43921 30619 43927
rect 23256 43862 24348 43890
rect 28000 43862 28212 43890
rect 23256 43850 23262 43862
rect 17402 43782 17408 43834
rect 17460 43782 17466 43834
rect 17954 43782 17960 43834
rect 18012 43822 18018 43834
rect 18693 43825 18751 43831
rect 18693 43822 18705 43825
rect 18012 43794 18705 43822
rect 18012 43782 18018 43794
rect 18693 43791 18705 43794
rect 18739 43791 18751 43825
rect 18693 43785 18751 43791
rect 19702 43782 19708 43834
rect 19760 43822 19766 43834
rect 21634 43822 21640 43834
rect 19760 43794 20116 43822
rect 19760 43782 19766 43794
rect 17586 43729 17592 43781
rect 17644 43729 17650 43781
rect 17862 43729 17868 43781
rect 17920 43729 17926 43781
rect 19337 43757 19395 43763
rect 19337 43723 19349 43757
rect 19383 43754 19395 43757
rect 19383 43726 19564 43754
rect 19383 43723 19395 43726
rect 19337 43717 19395 43723
rect 15764 43658 16891 43686
rect 15657 43649 15715 43655
rect 18782 43646 18788 43698
rect 18840 43686 18846 43698
rect 19429 43689 19487 43695
rect 19429 43686 19441 43689
rect 18840 43658 19441 43686
rect 18840 43646 18846 43658
rect 19429 43655 19441 43658
rect 19475 43655 19487 43689
rect 19536 43686 19564 43726
rect 19610 43714 19616 43766
rect 19668 43714 19674 43766
rect 19886 43714 19892 43766
rect 19944 43714 19950 43766
rect 20088 43763 20116 43794
rect 21100 43794 21640 43822
rect 20073 43757 20131 43763
rect 20073 43723 20085 43757
rect 20119 43723 20131 43757
rect 20073 43717 20131 43723
rect 20340 43757 20398 43763
rect 20340 43723 20352 43757
rect 20386 43754 20398 43757
rect 21100 43754 21128 43794
rect 21634 43782 21640 43794
rect 21692 43782 21698 43834
rect 22922 43782 22928 43834
rect 22980 43822 22986 43834
rect 24320 43822 24348 43862
rect 28184 43831 28212 43862
rect 28169 43825 28227 43831
rect 22980 43794 23980 43822
rect 24320 43794 24440 43822
rect 22980 43782 22986 43794
rect 23952 43782 23980 43794
rect 23952 43775 24072 43782
rect 23952 43769 24087 43775
rect 20386 43726 21128 43754
rect 20386 43723 20398 43726
rect 20340 43717 20398 43723
rect 19797 43689 19855 43695
rect 19797 43686 19809 43689
rect 19536 43658 19809 43686
rect 19429 43649 19487 43655
rect 19797 43655 19809 43658
rect 19843 43655 19855 43689
rect 20088 43686 20116 43717
rect 22646 43714 22652 43766
rect 22704 43763 22710 43766
rect 22704 43754 22716 43763
rect 22704 43726 22749 43754
rect 22704 43717 22716 43726
rect 22704 43714 22710 43717
rect 23382 43714 23388 43766
rect 23440 43714 23446 43766
rect 23477 43757 23535 43763
rect 23477 43723 23489 43757
rect 23523 43723 23535 43757
rect 23952 43754 24041 43769
rect 24029 43735 24041 43754
rect 24075 43754 24087 43769
rect 24305 43757 24363 43763
rect 24305 43754 24317 43757
rect 24075 43735 24317 43754
rect 24029 43729 24317 43735
rect 24044 43726 24317 43729
rect 23477 43717 23535 43723
rect 24305 43723 24317 43726
rect 24351 43723 24363 43757
rect 24412 43754 24440 43794
rect 28169 43791 28181 43825
rect 28215 43791 28227 43825
rect 28169 43785 28227 43791
rect 31110 43782 31116 43834
rect 31168 43782 31174 43834
rect 24578 43763 24584 43766
rect 24550 43757 24584 43763
rect 24550 43754 24562 43757
rect 24412 43726 24562 43754
rect 24305 43717 24363 43723
rect 24550 43723 24562 43726
rect 24550 43717 24584 43723
rect 22922 43686 22928 43698
rect 20088 43658 22928 43686
rect 19797 43649 19855 43655
rect 22922 43646 22928 43658
rect 22980 43646 22986 43698
rect 23014 43646 23020 43698
rect 23072 43646 23078 43698
rect 23198 43646 23204 43698
rect 23256 43686 23262 43698
rect 23492 43686 23520 43717
rect 23256 43658 23520 43686
rect 23256 43646 23262 43658
rect 23566 43646 23572 43698
rect 23624 43686 23630 43698
rect 23937 43689 23995 43695
rect 23937 43686 23949 43689
rect 23624 43658 23949 43686
rect 23624 43646 23630 43658
rect 23937 43655 23949 43658
rect 23983 43655 23995 43689
rect 24320 43686 24348 43717
rect 24578 43714 24584 43717
rect 24636 43714 24642 43766
rect 26878 43763 26884 43766
rect 26605 43757 26663 43763
rect 26605 43754 26617 43757
rect 24679 43726 26617 43754
rect 24394 43686 24400 43698
rect 24320 43658 24400 43686
rect 23937 43649 23995 43655
rect 24394 43646 24400 43658
rect 24452 43686 24458 43698
rect 24679 43686 24707 43726
rect 26605 43723 26617 43726
rect 26651 43723 26663 43757
rect 26605 43717 26663 43723
rect 26872 43717 26884 43763
rect 24452 43658 24707 43686
rect 24452 43646 24458 43658
rect 25498 43646 25504 43698
rect 25556 43686 25562 43698
rect 25685 43689 25743 43695
rect 25685 43686 25697 43689
rect 25556 43658 25697 43686
rect 25556 43646 25562 43658
rect 25685 43655 25697 43658
rect 25731 43655 25743 43689
rect 26620 43686 26648 43717
rect 26878 43714 26884 43717
rect 26936 43714 26942 43766
rect 28994 43754 29000 43766
rect 26988 43726 29000 43754
rect 26988 43686 27016 43726
rect 28994 43714 29000 43726
rect 29052 43714 29058 43766
rect 29270 43763 29276 43766
rect 29264 43717 29276 43763
rect 29270 43714 29276 43717
rect 29328 43714 29334 43766
rect 26620 43658 27016 43686
rect 25685 43649 25743 43655
rect 27982 43646 27988 43698
rect 28040 43646 28046 43698
rect 28350 43646 28356 43698
rect 28408 43646 28414 43698
rect 28445 43689 28503 43695
rect 28445 43655 28457 43689
rect 28491 43686 28503 43689
rect 28626 43686 28632 43698
rect 28491 43658 28632 43686
rect 28491 43655 28503 43658
rect 28445 43649 28503 43655
rect 28626 43646 28632 43658
rect 28684 43646 28690 43698
rect 28813 43689 28871 43695
rect 28813 43655 28825 43689
rect 28859 43686 28871 43689
rect 29362 43686 29368 43698
rect 28859 43658 29368 43686
rect 28859 43655 28871 43658
rect 28813 43649 28871 43655
rect 29362 43646 29368 43658
rect 29420 43646 29426 43698
rect 552 43546 31808 43568
rect 552 43494 8172 43546
rect 8224 43494 8236 43546
rect 8288 43494 8300 43546
rect 8352 43494 8364 43546
rect 8416 43494 8428 43546
rect 8480 43494 15946 43546
rect 15998 43494 16010 43546
rect 16062 43494 16074 43546
rect 16126 43494 16138 43546
rect 16190 43494 16202 43546
rect 16254 43494 23720 43546
rect 23772 43494 23784 43546
rect 23836 43494 23848 43546
rect 23900 43494 23912 43546
rect 23964 43494 23976 43546
rect 24028 43494 31494 43546
rect 31546 43494 31558 43546
rect 31610 43494 31622 43546
rect 31674 43494 31686 43546
rect 31738 43494 31750 43546
rect 31802 43494 31808 43546
rect 552 43472 31808 43494
rect 14182 43374 14188 43426
rect 14240 43374 14246 43426
rect 14461 43417 14519 43423
rect 14461 43414 14473 43417
rect 14292 43386 14473 43414
rect 13170 43306 13176 43358
rect 13228 43346 13234 43358
rect 14292 43346 14320 43386
rect 14461 43383 14473 43386
rect 14507 43414 14519 43417
rect 19242 43414 19248 43426
rect 14507 43386 15056 43414
rect 14507 43383 14519 43386
rect 14461 43377 14519 43383
rect 13228 43318 14320 43346
rect 13228 43306 13234 43318
rect 15028 43307 15056 43386
rect 15756 43386 19248 43414
rect 15013 43301 15071 43307
rect 13078 43238 13084 43290
rect 13136 43238 13142 43290
rect 13262 43238 13268 43290
rect 13320 43278 13326 43290
rect 14366 43287 14372 43290
rect 14344 43281 14372 43287
rect 14344 43278 14356 43281
rect 13320 43250 14356 43278
rect 13320 43238 13326 43250
rect 14344 43247 14356 43250
rect 14344 43241 14372 43247
rect 14366 43238 14372 43241
rect 14424 43238 14430 43290
rect 14829 43281 14887 43287
rect 14829 43247 14841 43281
rect 14875 43278 14887 43281
rect 14918 43278 14924 43290
rect 14875 43250 14924 43278
rect 14875 43247 14887 43250
rect 14829 43241 14887 43247
rect 14918 43238 14924 43250
rect 14976 43238 14982 43290
rect 15013 43267 15025 43301
rect 15059 43267 15071 43301
rect 15756 43295 15784 43386
rect 19242 43374 19248 43386
rect 19300 43374 19306 43426
rect 19334 43374 19340 43426
rect 19392 43374 19398 43426
rect 22646 43414 22652 43426
rect 16390 43355 16396 43358
rect 16384 43346 16396 43355
rect 16351 43318 16396 43346
rect 16384 43309 16396 43318
rect 16390 43306 16396 43309
rect 16448 43306 16454 43358
rect 18782 43306 18788 43358
rect 18840 43355 18846 43358
rect 18840 43346 18852 43355
rect 19352 43346 19380 43374
rect 18840 43318 18885 43346
rect 19076 43318 19380 43346
rect 19610 43340 19616 43392
rect 19668 43340 19674 43392
rect 20824 43386 22652 43414
rect 20824 43332 20852 43386
rect 22646 43374 22652 43386
rect 22704 43374 22710 43426
rect 22922 43374 22928 43426
rect 22980 43374 22986 43426
rect 23382 43374 23388 43426
rect 23440 43414 23446 43426
rect 25961 43417 26019 43423
rect 23440 43386 25912 43414
rect 23440 43374 23446 43386
rect 18840 43309 18852 43318
rect 18840 43306 18846 43309
rect 15013 43261 15071 43267
rect 15378 43238 15384 43290
rect 15436 43278 15442 43290
rect 15741 43289 15799 43295
rect 15741 43278 15753 43289
rect 15436 43255 15753 43278
rect 15787 43255 15799 43289
rect 19076 43287 19104 43318
rect 23198 43306 23204 43358
rect 23256 43346 23262 43358
rect 23814 43349 23872 43355
rect 23814 43346 23826 43349
rect 23256 43318 23826 43346
rect 23256 43306 23262 43318
rect 23814 43315 23826 43318
rect 23860 43315 23872 43349
rect 23814 43309 23872 43315
rect 23934 43306 23940 43358
rect 23992 43346 23998 43358
rect 23992 43318 24624 43346
rect 23992 43306 23998 43318
rect 15436 43250 15799 43255
rect 15436 43238 15442 43250
rect 15741 43249 15799 43250
rect 15841 43281 15899 43287
rect 15841 43247 15853 43281
rect 15887 43278 15899 43281
rect 16117 43281 16175 43287
rect 16117 43278 16129 43281
rect 15887 43250 16129 43278
rect 15887 43247 15899 43250
rect 15841 43241 15899 43247
rect 16117 43247 16129 43250
rect 16163 43247 16175 43281
rect 16117 43241 16175 43247
rect 19061 43281 19119 43287
rect 19061 43247 19073 43281
rect 19107 43247 19119 43281
rect 19061 43241 19119 43247
rect 19242 43238 19248 43290
rect 19300 43278 19306 43290
rect 19337 43281 19395 43287
rect 19337 43278 19349 43281
rect 19300 43250 19349 43278
rect 19300 43238 19306 43250
rect 19337 43247 19349 43250
rect 19383 43247 19395 43281
rect 19337 43241 19395 43247
rect 21450 43238 21456 43290
rect 21508 43238 21514 43290
rect 23566 43238 23572 43290
rect 23624 43238 23630 43290
rect 24596 43278 24624 43318
rect 24670 43306 24676 43358
rect 24728 43346 24734 43358
rect 25133 43349 25191 43355
rect 25133 43346 25145 43349
rect 24728 43318 25145 43346
rect 24728 43306 24734 43318
rect 25133 43315 25145 43318
rect 25179 43315 25191 43349
rect 25133 43309 25191 43315
rect 25498 43306 25504 43358
rect 25556 43306 25562 43358
rect 25884 43346 25912 43386
rect 25961 43383 25973 43417
rect 26007 43414 26019 43417
rect 26602 43414 26608 43426
rect 26007 43386 26608 43414
rect 26007 43383 26019 43386
rect 25961 43377 26019 43383
rect 26602 43374 26608 43386
rect 26660 43374 26666 43426
rect 26878 43374 26884 43426
rect 26936 43374 26942 43426
rect 28350 43374 28356 43426
rect 28408 43414 28414 43426
rect 28905 43417 28963 43423
rect 28905 43414 28917 43417
rect 28408 43386 28917 43414
rect 28408 43374 28414 43386
rect 28905 43383 28917 43386
rect 28951 43383 28963 43417
rect 28905 43377 28963 43383
rect 29181 43417 29239 43423
rect 29181 43383 29193 43417
rect 29227 43383 29239 43417
rect 29181 43377 29239 43383
rect 27982 43346 27988 43358
rect 25884 43318 27988 43346
rect 27982 43306 27988 43318
rect 28040 43306 28046 43358
rect 28568 43349 28626 43355
rect 28568 43315 28580 43349
rect 28614 43346 28626 43349
rect 29196 43346 29224 43377
rect 29546 43374 29552 43426
rect 29604 43414 29610 43426
rect 29604 43386 30604 43414
rect 29604 43374 29610 43386
rect 28614 43318 29224 43346
rect 29724 43349 29782 43355
rect 28614 43315 28626 43318
rect 28568 43309 28626 43315
rect 29724 43315 29736 43349
rect 29770 43346 29782 43349
rect 30466 43346 30472 43358
rect 29770 43318 30472 43346
rect 29770 43315 29782 43318
rect 29724 43309 29782 43315
rect 30466 43306 30472 43318
rect 30524 43306 30530 43358
rect 24596 43250 24992 43278
rect 11330 43170 11336 43222
rect 11388 43170 11394 43222
rect 12618 43170 12624 43222
rect 12676 43210 12682 43222
rect 13449 43213 13507 43219
rect 13449 43210 13461 43213
rect 12676 43182 13461 43210
rect 12676 43170 12682 43182
rect 13449 43179 13461 43182
rect 13495 43179 13507 43213
rect 13449 43173 13507 43179
rect 13538 43170 13544 43222
rect 13596 43210 13602 43222
rect 14553 43213 14611 43219
rect 14553 43210 14565 43213
rect 13596 43182 14565 43210
rect 13596 43170 13602 43182
rect 14553 43179 14565 43182
rect 14599 43210 14611 43213
rect 15286 43210 15292 43222
rect 14599 43182 15292 43210
rect 14599 43179 14611 43182
rect 14553 43173 14611 43179
rect 15286 43170 15292 43182
rect 15344 43170 15350 43222
rect 17310 43170 17316 43222
rect 17368 43210 17374 43222
rect 17681 43213 17739 43219
rect 17681 43210 17693 43213
rect 17368 43182 17693 43210
rect 17368 43170 17374 43182
rect 17681 43179 17693 43182
rect 17727 43210 17739 43213
rect 17954 43210 17960 43222
rect 17727 43182 17960 43210
rect 17727 43179 17739 43182
rect 17681 43173 17739 43179
rect 17954 43170 17960 43182
rect 18012 43170 18018 43222
rect 24964 43219 24992 43250
rect 25222 43246 25228 43298
rect 25280 43246 25286 43298
rect 25424 43250 26464 43278
rect 24949 43213 25007 43219
rect 24949 43179 24961 43213
rect 24995 43179 25007 43213
rect 24949 43173 25007 43179
rect 11790 43102 11796 43154
rect 11848 43142 11854 43154
rect 15194 43142 15200 43154
rect 11848 43114 15200 43142
rect 11848 43102 11854 43114
rect 15194 43102 15200 43114
rect 15252 43142 15258 43154
rect 16114 43142 16120 43154
rect 15252 43114 16120 43142
rect 15252 43102 15258 43114
rect 16114 43102 16120 43114
rect 16172 43102 16178 43154
rect 17034 43102 17040 43154
rect 17092 43142 17098 43154
rect 17497 43145 17555 43151
rect 17497 43142 17509 43145
rect 17092 43114 17509 43142
rect 17092 43102 17098 43114
rect 17497 43111 17509 43114
rect 17543 43111 17555 43145
rect 17497 43105 17555 43111
rect 21085 43145 21143 43151
rect 21085 43111 21097 43145
rect 21131 43142 21143 43145
rect 22554 43142 22560 43154
rect 21131 43114 22560 43142
rect 21131 43111 21143 43114
rect 21085 43105 21143 43111
rect 22554 43102 22560 43114
rect 22612 43102 22618 43154
rect 24964 43142 24992 43173
rect 25038 43170 25044 43222
rect 25096 43210 25102 43222
rect 25424 43210 25452 43250
rect 25096 43182 25452 43210
rect 25096 43170 25102 43182
rect 25501 43179 25559 43185
rect 25501 43145 25513 43179
rect 25547 43145 25559 43179
rect 26050 43170 26056 43222
rect 26108 43170 26114 43222
rect 26234 43170 26240 43222
rect 26292 43170 26298 43222
rect 26436 43210 26464 43250
rect 26510 43238 26516 43290
rect 26568 43278 26574 43290
rect 26605 43281 26663 43287
rect 26605 43278 26617 43281
rect 26568 43250 26617 43278
rect 26568 43238 26574 43250
rect 26605 43247 26617 43250
rect 26651 43247 26663 43281
rect 26605 43241 26663 43247
rect 27062 43238 27068 43290
rect 27120 43238 27126 43290
rect 28813 43281 28871 43287
rect 28813 43247 28825 43281
rect 28859 43247 28871 43281
rect 28813 43241 28871 43247
rect 27430 43210 27436 43222
rect 26436 43182 27436 43210
rect 27430 43170 27436 43182
rect 27488 43170 27494 43222
rect 28828 43210 28856 43241
rect 28902 43238 28908 43290
rect 28960 43278 28966 43290
rect 29089 43281 29147 43287
rect 29089 43278 29101 43281
rect 28960 43250 29101 43278
rect 28960 43238 28966 43250
rect 29089 43247 29101 43250
rect 29135 43247 29147 43281
rect 29089 43241 29147 43247
rect 29362 43238 29368 43290
rect 29420 43238 29426 43290
rect 29457 43281 29515 43287
rect 29457 43247 29469 43281
rect 29503 43247 29515 43281
rect 30576 43278 30604 43386
rect 30834 43374 30840 43426
rect 30892 43414 30898 43426
rect 30929 43417 30987 43423
rect 30929 43414 30941 43417
rect 30892 43386 30941 43414
rect 30892 43374 30898 43386
rect 30929 43383 30941 43386
rect 30975 43383 30987 43417
rect 30929 43377 30987 43383
rect 31113 43281 31171 43287
rect 31113 43278 31125 43281
rect 30576 43250 31125 43278
rect 29457 43241 29515 43247
rect 31113 43247 31125 43250
rect 31159 43247 31171 43281
rect 31113 43241 31171 43247
rect 28994 43210 29000 43222
rect 28828 43182 29000 43210
rect 28994 43170 29000 43182
rect 29052 43210 29058 43222
rect 29472 43210 29500 43241
rect 29052 43182 29500 43210
rect 29052 43170 29058 43182
rect 25501 43142 25559 43145
rect 24964 43139 25559 43142
rect 24964 43114 25544 43139
rect 26418 43102 26424 43154
rect 26476 43102 26482 43154
rect 30837 43145 30895 43151
rect 30837 43111 30849 43145
rect 30883 43142 30895 43145
rect 31110 43142 31116 43154
rect 30883 43114 31116 43142
rect 30883 43111 30895 43114
rect 30837 43105 30895 43111
rect 31110 43102 31116 43114
rect 31168 43102 31174 43154
rect 200 43002 31648 43024
rect 200 42950 206 43002
rect 514 42950 4285 43002
rect 4337 42950 4349 43002
rect 4401 42950 4413 43002
rect 4465 42950 4477 43002
rect 4529 42950 4541 43002
rect 4593 42950 12059 43002
rect 12111 42950 12123 43002
rect 12175 42950 12187 43002
rect 12239 42950 12251 43002
rect 12303 42950 12315 43002
rect 12367 42950 19833 43002
rect 19885 42950 19897 43002
rect 19949 42950 19961 43002
rect 20013 42950 20025 43002
rect 20077 42950 20089 43002
rect 20141 42950 27607 43002
rect 27659 42950 27671 43002
rect 27723 42950 27735 43002
rect 27787 42950 27799 43002
rect 27851 42950 27863 43002
rect 27915 42950 31648 43002
rect 200 42928 31648 42950
rect 11146 42830 11152 42882
rect 11204 42830 11210 42882
rect 11701 42873 11759 42879
rect 11701 42839 11713 42873
rect 11747 42870 11759 42873
rect 12434 42870 12440 42882
rect 11747 42842 12440 42870
rect 11747 42839 11759 42842
rect 11701 42833 11759 42839
rect 12434 42830 12440 42842
rect 12492 42830 12498 42882
rect 13078 42830 13084 42882
rect 13136 42870 13142 42882
rect 16853 42873 16911 42879
rect 16853 42870 16865 42873
rect 13136 42842 16865 42870
rect 13136 42830 13142 42842
rect 16853 42839 16865 42842
rect 16899 42870 16911 42873
rect 21450 42870 21456 42882
rect 16899 42842 21456 42870
rect 16899 42839 16911 42842
rect 16853 42833 16911 42839
rect 21450 42830 21456 42842
rect 21508 42830 21514 42882
rect 21818 42830 21824 42882
rect 21876 42870 21882 42882
rect 23385 42873 23443 42879
rect 23385 42870 23397 42873
rect 21876 42842 23397 42870
rect 21876 42830 21882 42842
rect 23385 42839 23397 42842
rect 23431 42839 23443 42873
rect 26418 42870 26424 42882
rect 23385 42833 23443 42839
rect 25516 42842 26424 42870
rect 12618 42762 12624 42814
rect 12676 42802 12682 42814
rect 12713 42805 12771 42811
rect 12713 42802 12725 42805
rect 12676 42774 12725 42802
rect 12676 42762 12682 42774
rect 12713 42771 12725 42774
rect 12759 42771 12771 42805
rect 12713 42765 12771 42771
rect 13354 42762 13360 42814
rect 13412 42802 13418 42814
rect 13412 42774 14780 42802
rect 13412 42762 13418 42774
rect 11977 42737 12035 42743
rect 11977 42734 11989 42737
rect 11256 42706 11989 42734
rect 11256 42675 11284 42706
rect 11977 42703 11989 42706
rect 12023 42703 12035 42737
rect 11977 42697 12035 42703
rect 12253 42737 12311 42743
rect 12253 42703 12265 42737
rect 12299 42734 12311 42737
rect 13372 42734 13400 42762
rect 14752 42743 14780 42774
rect 15197 42771 15255 42777
rect 12299 42706 13400 42734
rect 14737 42737 14795 42743
rect 12299 42703 12311 42706
rect 12253 42697 12311 42703
rect 14737 42703 14749 42737
rect 14783 42734 14795 42737
rect 14918 42734 14924 42746
rect 14783 42706 14924 42734
rect 14783 42703 14795 42706
rect 14737 42697 14795 42703
rect 14918 42694 14924 42706
rect 14976 42694 14982 42746
rect 15010 42694 15016 42746
rect 15068 42734 15074 42746
rect 15197 42737 15209 42771
rect 15243 42737 15255 42771
rect 15378 42762 15384 42814
rect 15436 42802 15442 42814
rect 24029 42805 24087 42811
rect 15436 42774 15884 42802
rect 15436 42762 15442 42774
rect 15197 42734 15255 42737
rect 15068 42731 15255 42734
rect 15068 42706 15240 42731
rect 15068 42694 15074 42706
rect 11241 42669 11299 42675
rect 11241 42635 11253 42669
rect 11287 42635 11299 42669
rect 11241 42629 11299 42635
rect 11793 42669 11851 42675
rect 11793 42635 11805 42669
rect 11839 42666 11851 42669
rect 12526 42666 12532 42678
rect 11839 42638 12532 42666
rect 11839 42635 11851 42638
rect 11793 42629 11851 42635
rect 12526 42626 12532 42638
rect 12584 42626 12590 42678
rect 12713 42635 12771 42641
rect 12158 42558 12164 42610
rect 12216 42558 12222 42610
rect 12342 42558 12348 42610
rect 12400 42598 12406 42610
rect 12713 42601 12725 42635
rect 12759 42601 12771 42635
rect 12986 42626 12992 42678
rect 13044 42626 13050 42678
rect 13078 42626 13084 42678
rect 13136 42666 13142 42678
rect 13357 42669 13415 42675
rect 13357 42666 13369 42669
rect 13136 42638 13369 42666
rect 13136 42626 13142 42638
rect 13357 42635 13369 42638
rect 13403 42635 13415 42669
rect 13446 42641 13452 42693
rect 13504 42681 13510 42693
rect 15856 42690 15884 42774
rect 19536 42774 23888 42802
rect 16942 42694 16948 42746
rect 17000 42734 17006 42746
rect 17000 42706 18460 42734
rect 17000 42694 17006 42706
rect 13679 42684 13737 42690
rect 13679 42681 13691 42684
rect 13504 42653 13691 42681
rect 13504 42641 13510 42653
rect 13679 42650 13691 42653
rect 13725 42650 13737 42684
rect 13679 42644 13737 42650
rect 14277 42684 14335 42690
rect 14277 42650 14289 42684
rect 14323 42666 14335 42684
rect 15841 42684 15899 42690
rect 15194 42666 15200 42678
rect 14323 42650 15200 42666
rect 14277 42644 15200 42650
rect 14292 42638 15200 42644
rect 13357 42629 13415 42635
rect 15194 42626 15200 42638
rect 15252 42626 15258 42678
rect 15286 42626 15292 42678
rect 15344 42666 15350 42678
rect 15565 42669 15623 42675
rect 15344 42638 15516 42666
rect 15344 42626 15350 42638
rect 12713 42598 12771 42601
rect 13538 42598 13544 42610
rect 12400 42570 13544 42598
rect 12400 42558 12406 42570
rect 13538 42558 13544 42570
rect 13596 42558 13602 42610
rect 14182 42558 14188 42610
rect 14240 42558 14246 42610
rect 14921 42601 14979 42607
rect 14921 42567 14933 42601
rect 14967 42598 14979 42601
rect 15378 42598 15384 42610
rect 14967 42570 15384 42598
rect 14967 42567 14979 42570
rect 14921 42561 14979 42567
rect 15378 42558 15384 42570
rect 15436 42558 15442 42610
rect 15488 42598 15516 42638
rect 15565 42635 15577 42669
rect 15611 42666 15623 42669
rect 15654 42666 15660 42678
rect 15611 42638 15660 42666
rect 15611 42635 15623 42638
rect 15565 42629 15623 42635
rect 15654 42626 15660 42638
rect 15712 42626 15718 42678
rect 15841 42650 15853 42684
rect 15887 42650 15899 42684
rect 15841 42644 15899 42650
rect 16298 42641 16304 42693
rect 16356 42641 16362 42693
rect 18432 42675 18460 42706
rect 18141 42669 18199 42675
rect 18141 42635 18153 42669
rect 18187 42666 18199 42669
rect 18417 42669 18475 42675
rect 18187 42638 18368 42666
rect 18187 42635 18199 42638
rect 18141 42629 18199 42635
rect 17310 42598 17316 42610
rect 15488 42570 17316 42598
rect 17310 42558 17316 42570
rect 17368 42558 17374 42610
rect 18230 42558 18236 42610
rect 18288 42558 18294 42610
rect 18340 42598 18368 42638
rect 18417 42635 18429 42669
rect 18463 42635 18475 42669
rect 18417 42629 18475 42635
rect 19536 42598 19564 42774
rect 19610 42694 19616 42746
rect 19668 42734 19674 42746
rect 20898 42734 20904 42746
rect 19668 42706 20904 42734
rect 19668 42694 19674 42706
rect 20898 42694 20904 42706
rect 20956 42694 20962 42746
rect 20993 42737 21051 42743
rect 20993 42703 21005 42737
rect 21039 42703 21051 42737
rect 20993 42697 21051 42703
rect 21008 42666 21036 42697
rect 21082 42694 21088 42746
rect 21140 42734 21146 42746
rect 21269 42737 21327 42743
rect 21269 42734 21281 42737
rect 21140 42706 21281 42734
rect 21140 42694 21146 42706
rect 21269 42703 21281 42706
rect 21315 42703 21327 42737
rect 21269 42697 21327 42703
rect 21818 42694 21824 42746
rect 21876 42694 21882 42746
rect 22554 42694 22560 42746
rect 22612 42694 22618 42746
rect 23109 42737 23167 42743
rect 23109 42703 23121 42737
rect 23155 42734 23167 42737
rect 23474 42734 23480 42746
rect 23155 42706 23480 42734
rect 23155 42703 23167 42706
rect 23109 42697 23167 42703
rect 23474 42694 23480 42706
rect 23532 42694 23538 42746
rect 23860 42734 23888 42774
rect 24029 42771 24041 42805
rect 24075 42802 24087 42805
rect 24118 42802 24124 42814
rect 24075 42774 24124 42802
rect 24075 42771 24087 42774
rect 24029 42765 24087 42771
rect 24118 42762 24124 42774
rect 24176 42762 24182 42814
rect 23584 42706 23796 42734
rect 23860 42706 24256 42734
rect 22370 42666 22376 42678
rect 21008 42638 22376 42666
rect 22370 42626 22376 42638
rect 22428 42666 22434 42678
rect 22428 42638 23152 42666
rect 22428 42626 22434 42638
rect 18340 42570 19564 42598
rect 19886 42558 19892 42610
rect 19944 42598 19950 42610
rect 20441 42601 20499 42607
rect 20441 42598 20453 42601
rect 19944 42570 20453 42598
rect 19944 42558 19950 42570
rect 20441 42567 20453 42570
rect 20487 42567 20499 42601
rect 20441 42561 20499 42567
rect 20806 42558 20812 42610
rect 20864 42558 20870 42610
rect 20901 42601 20959 42607
rect 20901 42567 20913 42601
rect 20947 42598 20959 42601
rect 21174 42598 21180 42610
rect 20947 42570 21180 42598
rect 20947 42567 20959 42570
rect 20901 42561 20959 42567
rect 21174 42558 21180 42570
rect 21232 42558 21238 42610
rect 21450 42558 21456 42610
rect 21508 42598 21514 42610
rect 22005 42601 22063 42607
rect 22005 42598 22017 42601
rect 21508 42570 22017 42598
rect 21508 42558 21514 42570
rect 22005 42567 22017 42570
rect 22051 42567 22063 42601
rect 22005 42561 22063 42567
rect 22738 42558 22744 42610
rect 22796 42598 22802 42610
rect 23014 42598 23020 42610
rect 22796 42570 23020 42598
rect 22796 42558 22802 42570
rect 23014 42558 23020 42570
rect 23072 42558 23078 42610
rect 23124 42598 23152 42638
rect 23198 42626 23204 42678
rect 23256 42626 23262 42678
rect 23584 42666 23612 42706
rect 23308 42638 23612 42666
rect 23661 42669 23719 42675
rect 23308 42598 23336 42638
rect 23661 42635 23673 42669
rect 23707 42635 23719 42669
rect 23768 42666 23796 42706
rect 23934 42666 23940 42678
rect 23768 42638 23940 42666
rect 23661 42629 23719 42635
rect 23124 42570 23336 42598
rect 23474 42558 23480 42610
rect 23532 42558 23538 42610
rect 23676 42598 23704 42629
rect 23934 42626 23940 42638
rect 23992 42626 23998 42678
rect 23845 42601 23903 42607
rect 23845 42598 23857 42601
rect 23676 42570 23857 42598
rect 23845 42567 23857 42570
rect 23891 42567 23903 42601
rect 24228 42598 24256 42706
rect 24394 42694 24400 42746
rect 24452 42694 24458 42746
rect 24305 42669 24363 42675
rect 24305 42635 24317 42669
rect 24351 42666 24363 42669
rect 24486 42666 24492 42678
rect 24351 42638 24492 42666
rect 24351 42635 24363 42638
rect 24305 42629 24363 42635
rect 24486 42626 24492 42638
rect 24544 42626 24550 42678
rect 24664 42669 24722 42675
rect 24664 42635 24676 42669
rect 24710 42666 24722 42669
rect 25516 42666 25544 42842
rect 26418 42830 26424 42842
rect 26476 42830 26482 42882
rect 28626 42830 28632 42882
rect 28684 42830 28690 42882
rect 29178 42830 29184 42882
rect 29236 42830 29242 42882
rect 29270 42830 29276 42882
rect 29328 42830 29334 42882
rect 30466 42830 30472 42882
rect 30524 42830 30530 42882
rect 30926 42802 30932 42814
rect 24710 42638 25544 42666
rect 25700 42774 30932 42802
rect 24710 42635 24722 42638
rect 24664 42629 24722 42635
rect 25700 42598 25728 42774
rect 30926 42762 30932 42774
rect 30984 42762 30990 42814
rect 26421 42737 26479 42743
rect 26421 42734 26433 42737
rect 25792 42706 26433 42734
rect 25792 42607 25820 42706
rect 26421 42703 26433 42706
rect 26467 42703 26479 42737
rect 26421 42697 26479 42703
rect 27430 42694 27436 42746
rect 27488 42734 27494 42746
rect 27985 42737 28043 42743
rect 27985 42734 27997 42737
rect 27488 42706 27997 42734
rect 27488 42694 27494 42706
rect 27985 42703 27997 42706
rect 28031 42703 28043 42737
rect 27985 42697 28043 42703
rect 26050 42626 26056 42678
rect 26108 42666 26114 42678
rect 26605 42669 26663 42675
rect 26605 42666 26617 42669
rect 26108 42638 26617 42666
rect 26108 42626 26114 42638
rect 26605 42635 26617 42638
rect 26651 42635 26663 42669
rect 26605 42629 26663 42635
rect 26786 42626 26792 42678
rect 26844 42626 26850 42678
rect 28810 42626 28816 42678
rect 28868 42666 28874 42678
rect 28997 42669 29055 42675
rect 28997 42666 29009 42669
rect 28868 42638 29009 42666
rect 28868 42626 28874 42638
rect 28997 42635 29009 42638
rect 29043 42635 29055 42669
rect 28997 42629 29055 42635
rect 29454 42626 29460 42678
rect 29512 42626 29518 42678
rect 30558 42626 30564 42678
rect 30616 42666 30622 42678
rect 30653 42669 30711 42675
rect 30653 42666 30665 42669
rect 30616 42638 30665 42666
rect 30616 42626 30622 42638
rect 30653 42635 30665 42638
rect 30699 42635 30711 42669
rect 30653 42629 30711 42635
rect 24228 42570 25728 42598
rect 25777 42601 25835 42607
rect 23845 42561 23903 42567
rect 25777 42567 25789 42601
rect 25823 42567 25835 42601
rect 25777 42561 25835 42567
rect 25866 42558 25872 42610
rect 25924 42558 25930 42610
rect 552 42458 31808 42480
rect 552 42406 8172 42458
rect 8224 42406 8236 42458
rect 8288 42406 8300 42458
rect 8352 42406 8364 42458
rect 8416 42406 8428 42458
rect 8480 42406 15946 42458
rect 15998 42406 16010 42458
rect 16062 42406 16074 42458
rect 16126 42406 16138 42458
rect 16190 42406 16202 42458
rect 16254 42406 23720 42458
rect 23772 42406 23784 42458
rect 23836 42406 23848 42458
rect 23900 42406 23912 42458
rect 23964 42406 23976 42458
rect 24028 42406 31494 42458
rect 31546 42406 31558 42458
rect 31610 42406 31622 42458
rect 31674 42406 31686 42458
rect 31738 42406 31750 42458
rect 31802 42406 31808 42458
rect 552 42384 31808 42406
rect 11514 42286 11520 42338
rect 11572 42326 11578 42338
rect 12069 42329 12127 42335
rect 12069 42326 12081 42329
rect 11572 42298 12081 42326
rect 11572 42286 11578 42298
rect 12069 42295 12081 42298
rect 12115 42295 12127 42329
rect 12069 42289 12127 42295
rect 12342 42286 12348 42338
rect 12400 42286 12406 42338
rect 12894 42286 12900 42338
rect 12952 42326 12958 42338
rect 13173 42329 13231 42335
rect 13173 42326 13185 42329
rect 12952 42298 13185 42326
rect 12952 42286 12958 42298
rect 13173 42295 13185 42298
rect 13219 42326 13231 42329
rect 13446 42326 13452 42338
rect 13219 42298 13452 42326
rect 13219 42295 13231 42298
rect 13173 42289 13231 42295
rect 13446 42286 13452 42298
rect 13504 42286 13510 42338
rect 13538 42286 13544 42338
rect 13596 42286 13602 42338
rect 13814 42286 13820 42338
rect 13872 42326 13878 42338
rect 14274 42326 14280 42338
rect 13872 42298 14280 42326
rect 13872 42286 13878 42298
rect 14274 42286 14280 42298
rect 14332 42286 14338 42338
rect 14458 42286 14464 42338
rect 14516 42326 14522 42338
rect 14516 42298 16344 42326
rect 14516 42286 14522 42298
rect 2314 42218 2320 42270
rect 2372 42258 2378 42270
rect 2970 42261 3028 42267
rect 2970 42258 2982 42261
rect 2372 42230 2982 42258
rect 2372 42218 2378 42230
rect 2970 42227 2982 42230
rect 3016 42227 3028 42261
rect 3878 42258 3884 42270
rect 2970 42221 3028 42227
rect 3252 42230 3884 42258
rect 3252 42199 3280 42230
rect 3878 42218 3884 42230
rect 3936 42258 3942 42270
rect 11330 42258 11336 42270
rect 3936 42230 11336 42258
rect 3936 42218 3942 42230
rect 11330 42218 11336 42230
rect 11388 42218 11394 42270
rect 11793 42261 11851 42267
rect 11793 42227 11805 42261
rect 11839 42258 11851 42261
rect 12158 42258 12164 42270
rect 11839 42230 12164 42258
rect 11839 42227 11851 42230
rect 11793 42221 11851 42227
rect 12158 42218 12164 42230
rect 12216 42258 12222 42270
rect 12253 42261 12311 42267
rect 12253 42258 12265 42261
rect 12216 42230 12265 42258
rect 12216 42218 12222 42230
rect 12253 42227 12265 42230
rect 12299 42258 12311 42261
rect 12805 42261 12863 42267
rect 12299 42230 12731 42258
rect 12299 42227 12311 42230
rect 12253 42221 12311 42227
rect 3237 42193 3295 42199
rect 3237 42159 3249 42193
rect 3283 42159 3295 42193
rect 3237 42153 3295 42159
rect 3418 42150 3424 42202
rect 3476 42150 3482 42202
rect 12703 42198 12731 42230
rect 12805 42227 12817 42261
rect 12851 42258 12863 42261
rect 12851 42230 13400 42258
rect 12851 42227 12863 42230
rect 12805 42221 12863 42227
rect 13372 42202 13400 42230
rect 12703 42190 12756 42198
rect 12989 42193 13047 42199
rect 12989 42190 13001 42193
rect 12703 42170 13001 42190
rect 12728 42162 13001 42170
rect 12989 42159 13001 42162
rect 13035 42159 13047 42193
rect 12989 42153 13047 42159
rect 11425 42125 11483 42131
rect 11425 42091 11437 42125
rect 11471 42122 11483 42125
rect 12618 42122 12624 42134
rect 11471 42094 12624 42122
rect 11471 42091 11483 42094
rect 11425 42085 11483 42091
rect 12618 42082 12624 42094
rect 12676 42082 12682 42134
rect 13004 42122 13032 42153
rect 13354 42150 13360 42202
rect 13412 42190 13418 42202
rect 13556 42199 13584 42286
rect 13998 42218 14004 42270
rect 14056 42258 14062 42270
rect 14056 42230 14964 42258
rect 14056 42218 14062 42230
rect 14553 42227 14611 42230
rect 13468 42193 13526 42199
rect 13468 42190 13480 42193
rect 13412 42162 13480 42190
rect 13412 42150 13418 42162
rect 13468 42159 13480 42162
rect 13514 42159 13526 42193
rect 13556 42193 13624 42199
rect 13556 42162 13578 42193
rect 13468 42153 13526 42159
rect 13566 42159 13578 42162
rect 13612 42159 13624 42193
rect 13566 42153 13624 42159
rect 14093 42193 14151 42199
rect 14093 42159 14105 42193
rect 14139 42190 14151 42193
rect 14182 42190 14188 42202
rect 14139 42162 14188 42190
rect 14139 42159 14151 42162
rect 14093 42153 14151 42159
rect 14182 42150 14188 42162
rect 14240 42150 14246 42202
rect 14366 42150 14372 42202
rect 14424 42150 14430 42202
rect 14553 42193 14565 42227
rect 14599 42193 14611 42227
rect 14553 42187 14611 42193
rect 14936 42211 14964 42230
rect 15197 42214 15255 42220
rect 15197 42211 15209 42214
rect 14936 42202 15209 42211
rect 14936 42183 15108 42202
rect 15102 42150 15108 42183
rect 15160 42183 15209 42202
rect 15160 42150 15166 42183
rect 15197 42180 15209 42183
rect 15243 42180 15255 42214
rect 15197 42174 15255 42180
rect 15378 42171 15384 42223
rect 15436 42211 15442 42223
rect 15654 42211 15660 42223
rect 15436 42183 15660 42211
rect 15436 42171 15442 42183
rect 15654 42171 15660 42183
rect 15712 42171 15718 42223
rect 16316 42199 16344 42298
rect 16390 42286 16396 42338
rect 16448 42326 16454 42338
rect 22097 42329 22155 42335
rect 22097 42326 22109 42329
rect 16448 42298 20024 42326
rect 16448 42286 16454 42298
rect 19996 42292 20024 42298
rect 20180 42298 22109 42326
rect 20180 42292 20208 42298
rect 16301 42193 16359 42199
rect 16301 42159 16313 42193
rect 16347 42159 16359 42193
rect 16942 42166 16948 42218
rect 17000 42206 17006 42218
rect 17036 42209 17094 42215
rect 17036 42206 17048 42209
rect 17000 42178 17048 42206
rect 17000 42166 17006 42178
rect 17036 42175 17048 42178
rect 17082 42175 17094 42209
rect 17036 42169 17094 42175
rect 16301 42153 16359 42159
rect 17126 42150 17132 42202
rect 17184 42190 17190 42202
rect 17221 42193 17279 42199
rect 17221 42190 17233 42193
rect 17184 42162 17233 42190
rect 17184 42150 17190 42162
rect 17221 42159 17233 42162
rect 17267 42159 17279 42193
rect 17310 42174 17316 42226
rect 17368 42174 17374 42226
rect 17402 42218 17408 42270
rect 17460 42258 17466 42270
rect 19794 42258 19800 42270
rect 17460 42230 19800 42258
rect 17460 42218 17466 42230
rect 19794 42218 19800 42230
rect 19852 42218 19858 42270
rect 19996 42264 20208 42292
rect 22097 42295 22109 42298
rect 22143 42295 22155 42329
rect 22097 42289 22155 42295
rect 22738 42286 22744 42338
rect 22796 42286 22802 42338
rect 23290 42286 23296 42338
rect 23348 42326 23354 42338
rect 23385 42329 23443 42335
rect 23385 42326 23397 42329
rect 23348 42298 23397 42326
rect 23348 42286 23354 42298
rect 23385 42295 23397 42298
rect 23431 42295 23443 42329
rect 23385 42289 23443 42295
rect 24302 42286 24308 42338
rect 24360 42326 24366 42338
rect 25406 42326 25412 42338
rect 24360 42298 25412 42326
rect 24360 42286 24366 42298
rect 20073 42227 20131 42233
rect 20073 42224 20085 42227
rect 19613 42193 19671 42199
rect 19613 42190 19625 42193
rect 17221 42153 17279 42159
rect 17788 42162 19625 42190
rect 14384 42122 14412 42150
rect 1854 42014 1860 42066
rect 1912 42014 1918 42066
rect 4065 42057 4123 42063
rect 4065 42023 4077 42057
rect 4111 42054 4123 42057
rect 4154 42054 4160 42066
rect 4111 42026 4160 42054
rect 4111 42023 4123 42026
rect 4065 42017 4123 42023
rect 4154 42014 4160 42026
rect 4212 42014 4218 42066
rect 11790 41964 11796 42016
rect 11848 41964 11854 42016
rect 11974 42014 11980 42066
rect 12032 42014 12038 42066
rect 12710 42048 12716 42100
rect 12768 42088 12774 42100
rect 12805 42091 12863 42097
rect 13004 42094 14412 42122
rect 14737 42125 14795 42131
rect 12805 42088 12817 42091
rect 12768 42060 12817 42088
rect 12768 42048 12774 42060
rect 12805 42057 12817 42060
rect 12851 42057 12863 42091
rect 13832 42066 13860 42094
rect 14737 42091 14749 42125
rect 14783 42122 14795 42125
rect 15470 42122 15476 42134
rect 14783 42094 15476 42122
rect 14783 42091 14795 42094
rect 14737 42085 14795 42091
rect 15470 42082 15476 42094
rect 15528 42082 15534 42134
rect 15562 42082 15568 42134
rect 15620 42122 15626 42134
rect 15657 42125 15715 42131
rect 15657 42122 15669 42125
rect 15620 42094 15669 42122
rect 15620 42082 15626 42094
rect 15657 42091 15669 42094
rect 15703 42122 15715 42125
rect 16485 42125 16543 42131
rect 15703 42094 16436 42122
rect 15703 42091 15715 42094
rect 15657 42085 15715 42091
rect 12805 42054 12863 42057
rect 12986 42054 12992 42066
rect 12805 42051 12992 42054
rect 12820 42026 12992 42051
rect 12986 42014 12992 42026
rect 13044 42014 13050 42066
rect 13814 42014 13820 42066
rect 13872 42014 13878 42066
rect 14274 41964 14280 42016
rect 14332 41964 14338 42016
rect 14826 42014 14832 42066
rect 14884 42054 14890 42066
rect 16117 42057 16175 42063
rect 16117 42054 16129 42057
rect 14884 42026 16129 42054
rect 14884 42014 14890 42026
rect 16117 42023 16129 42026
rect 16163 42023 16175 42057
rect 16408 42054 16436 42094
rect 16485 42091 16497 42125
rect 16531 42122 16543 42125
rect 16574 42122 16580 42134
rect 16531 42094 16580 42122
rect 16531 42091 16543 42094
rect 16485 42085 16543 42091
rect 16574 42082 16580 42094
rect 16632 42082 16638 42134
rect 16850 42082 16856 42134
rect 16908 42082 16914 42134
rect 17788 42122 17816 42162
rect 19613 42159 19625 42162
rect 19659 42159 19671 42193
rect 19613 42153 19671 42159
rect 19886 42150 19892 42202
rect 19944 42190 19950 42202
rect 19996 42196 20085 42224
rect 19996 42190 20024 42196
rect 19944 42162 20024 42190
rect 20073 42193 20085 42196
rect 20119 42193 20131 42227
rect 20254 42218 20260 42270
rect 20312 42218 20318 42270
rect 20346 42218 20352 42270
rect 20404 42258 20410 42270
rect 20404 42230 20760 42258
rect 20404 42218 20410 42230
rect 20732 42199 20760 42230
rect 20073 42187 20131 42193
rect 20441 42193 20499 42199
rect 19944 42150 19950 42162
rect 20441 42159 20453 42193
rect 20487 42190 20499 42193
rect 20625 42193 20683 42199
rect 20625 42190 20637 42193
rect 20487 42162 20637 42190
rect 20487 42159 20499 42162
rect 20441 42153 20499 42159
rect 20625 42159 20637 42162
rect 20671 42159 20683 42193
rect 20625 42153 20683 42159
rect 20717 42193 20775 42199
rect 20717 42159 20729 42193
rect 20763 42159 20775 42193
rect 21450 42184 21456 42236
rect 21508 42184 21514 42236
rect 21634 42218 21640 42270
rect 21692 42218 21698 42270
rect 21739 42227 21797 42233
rect 21637 42193 21649 42218
rect 21683 42193 21695 42218
rect 21637 42187 21695 42193
rect 21739 42193 21751 42227
rect 21785 42224 21797 42227
rect 21910 42224 21916 42236
rect 21785 42196 21916 42224
rect 21785 42193 21797 42196
rect 21739 42187 21797 42193
rect 21910 42184 21916 42196
rect 21968 42184 21974 42236
rect 22278 42218 22284 42270
rect 22336 42218 22342 42270
rect 24578 42258 24584 42270
rect 23124 42230 24584 42258
rect 22370 42166 22376 42218
rect 22428 42166 22434 42218
rect 22462 42166 22468 42218
rect 22520 42206 22526 42218
rect 22557 42209 22615 42215
rect 22557 42206 22569 42209
rect 22520 42178 22569 42206
rect 22520 42166 22526 42178
rect 22557 42175 22569 42178
rect 22603 42175 22615 42209
rect 23124 42199 23152 42230
rect 24578 42218 24584 42230
rect 24636 42218 24642 42270
rect 24745 42227 24803 42233
rect 22557 42169 22615 42175
rect 23109 42193 23167 42199
rect 20717 42153 20775 42159
rect 23109 42159 23121 42193
rect 23155 42159 23167 42193
rect 23109 42153 23167 42159
rect 17144 42094 17816 42122
rect 17144 42054 17172 42094
rect 18046 42082 18052 42134
rect 18104 42122 18110 42134
rect 19242 42122 19248 42134
rect 18104 42094 19248 42122
rect 18104 42082 18110 42094
rect 19242 42082 19248 42094
rect 19300 42122 19306 42134
rect 19426 42122 19432 42134
rect 19300 42094 19432 42122
rect 19300 42082 19306 42094
rect 19426 42082 19432 42094
rect 19484 42082 19490 42134
rect 19797 42125 19855 42131
rect 19797 42091 19809 42125
rect 19843 42122 19855 42125
rect 20640 42122 20668 42153
rect 23198 42150 23204 42202
rect 23256 42150 23262 42202
rect 24210 42150 24216 42202
rect 24268 42190 24274 42202
rect 24489 42193 24547 42199
rect 24489 42190 24501 42193
rect 24268 42162 24501 42190
rect 24268 42150 24274 42162
rect 24489 42159 24501 42162
rect 24535 42159 24547 42193
rect 24745 42193 24757 42227
rect 24791 42224 24803 42227
rect 24872 42224 24900 42298
rect 25406 42286 25412 42298
rect 25464 42326 25470 42338
rect 25866 42326 25872 42338
rect 25464 42298 25872 42326
rect 25464 42286 25470 42298
rect 25866 42286 25872 42298
rect 25924 42286 25930 42338
rect 24791 42196 24900 42224
rect 24791 42193 24803 42196
rect 24745 42187 24803 42193
rect 26973 42193 27031 42199
rect 24489 42153 24547 42159
rect 26973 42159 26985 42193
rect 27019 42159 27031 42193
rect 26973 42153 27031 42159
rect 20806 42122 20812 42134
rect 19843 42094 20576 42122
rect 20640 42094 20812 42122
rect 19843 42091 19855 42094
rect 19797 42085 19855 42091
rect 16408 42026 17172 42054
rect 19889 42057 19947 42063
rect 16117 42017 16175 42023
rect 19889 42023 19901 42057
rect 19935 42054 19947 42057
rect 20070 42054 20076 42066
rect 19935 42026 20076 42054
rect 19935 42023 19947 42026
rect 19889 42017 19947 42023
rect 20070 42014 20076 42026
rect 20128 42014 20134 42066
rect 20548 42054 20576 42094
rect 20806 42082 20812 42094
rect 20864 42122 20870 42134
rect 21082 42122 21088 42134
rect 20864 42094 21088 42122
rect 20864 42082 20870 42094
rect 21082 42082 21088 42094
rect 21140 42082 21146 42134
rect 21269 42125 21327 42131
rect 21269 42091 21281 42125
rect 21315 42122 21327 42125
rect 21818 42122 21824 42134
rect 21315 42094 21824 42122
rect 21315 42091 21327 42094
rect 21269 42085 21327 42091
rect 21818 42082 21824 42094
rect 21876 42082 21882 42134
rect 22646 42122 22652 42134
rect 22388 42094 22652 42122
rect 20714 42054 20720 42066
rect 20548 42026 20720 42054
rect 20714 42014 20720 42026
rect 20772 42014 20778 42066
rect 20898 42014 20904 42066
rect 20956 42014 20962 42066
rect 21358 42014 21364 42066
rect 21416 42054 21422 42066
rect 21913 42057 21971 42063
rect 21913 42054 21925 42057
rect 21416 42026 21925 42054
rect 21416 42014 21422 42026
rect 21913 42023 21925 42026
rect 21959 42023 21971 42057
rect 21913 42017 21971 42023
rect 22131 42007 22189 42013
rect 22131 41973 22143 42007
rect 22177 42004 22189 42007
rect 22388 42004 22416 42094
rect 22646 42082 22652 42094
rect 22704 42082 22710 42134
rect 25869 42125 25927 42131
rect 25869 42091 25881 42125
rect 25915 42122 25927 42125
rect 26988 42122 27016 42153
rect 25915 42094 27016 42122
rect 25915 42091 25927 42094
rect 25869 42085 25927 42091
rect 22462 42014 22468 42066
rect 22520 42054 22526 42066
rect 22557 42057 22615 42063
rect 22557 42054 22569 42057
rect 22520 42026 22569 42054
rect 22520 42014 22526 42026
rect 22557 42023 22569 42026
rect 22603 42023 22615 42057
rect 22557 42017 22615 42023
rect 25682 42014 25688 42066
rect 25740 42054 25746 42066
rect 26421 42057 26479 42063
rect 26421 42054 26433 42057
rect 25740 42026 26433 42054
rect 25740 42014 25746 42026
rect 26421 42023 26433 42026
rect 26467 42023 26479 42057
rect 26421 42017 26479 42023
rect 22177 41976 22416 42004
rect 22177 41973 22189 41976
rect 22131 41967 22189 41973
rect 200 41914 31648 41936
rect 200 41862 206 41914
rect 514 41862 4285 41914
rect 4337 41862 4349 41914
rect 4401 41862 4413 41914
rect 4465 41862 4477 41914
rect 4529 41862 4541 41914
rect 4593 41862 12059 41914
rect 12111 41862 12123 41914
rect 12175 41862 12187 41914
rect 12239 41862 12251 41914
rect 12303 41862 12315 41914
rect 12367 41862 19833 41914
rect 19885 41862 19897 41914
rect 19949 41862 19961 41914
rect 20013 41862 20025 41914
rect 20077 41862 20089 41914
rect 20141 41862 27607 41914
rect 27659 41862 27671 41914
rect 27723 41862 27735 41914
rect 27787 41862 27799 41914
rect 27851 41862 27863 41914
rect 27915 41862 31648 41914
rect 200 41840 31648 41862
rect 12342 41742 12348 41794
rect 12400 41782 12406 41794
rect 14185 41785 14243 41791
rect 14185 41782 14197 41785
rect 12400 41754 14197 41782
rect 12400 41742 12406 41754
rect 14185 41751 14197 41754
rect 14231 41782 14243 41785
rect 14550 41782 14556 41794
rect 14231 41754 14556 41782
rect 14231 41751 14243 41754
rect 14185 41745 14243 41751
rect 14550 41742 14556 41754
rect 14608 41742 14614 41794
rect 16298 41782 16304 41794
rect 14936 41754 16304 41782
rect 6641 41717 6699 41723
rect 6641 41683 6653 41717
rect 6687 41714 6699 41717
rect 14936 41714 14964 41754
rect 16298 41742 16304 41754
rect 16356 41742 16362 41794
rect 16942 41782 16948 41794
rect 16408 41754 16948 41782
rect 6687 41686 14964 41714
rect 6687 41683 6699 41686
rect 6641 41677 6699 41683
rect 15010 41674 15016 41726
rect 15068 41714 15074 41726
rect 16408 41714 16436 41754
rect 16942 41742 16948 41754
rect 17000 41742 17006 41794
rect 17218 41742 17224 41794
rect 17276 41782 17282 41794
rect 17276 41754 19472 41782
rect 17276 41742 17282 41754
rect 15068 41689 16436 41714
rect 15068 41686 16451 41689
rect 15068 41674 15074 41686
rect 16393 41683 16451 41686
rect 1854 41606 1860 41658
rect 1912 41646 1918 41658
rect 2409 41649 2467 41655
rect 2409 41646 2421 41649
rect 1912 41618 2421 41646
rect 1912 41606 1918 41618
rect 2409 41615 2421 41618
rect 2455 41615 2467 41649
rect 2409 41609 2467 41615
rect 5258 41606 5264 41658
rect 5316 41646 5322 41658
rect 5997 41649 6055 41655
rect 5997 41646 6009 41649
rect 5316 41618 6009 41646
rect 5316 41606 5322 41618
rect 5997 41615 6009 41618
rect 6043 41615 6055 41649
rect 5997 41609 6055 41615
rect 13078 41606 13084 41658
rect 13136 41646 13142 41658
rect 13630 41646 13636 41658
rect 13136 41618 13636 41646
rect 13136 41606 13142 41618
rect 13630 41606 13636 41618
rect 13688 41606 13694 41658
rect 13725 41609 13783 41615
rect 12023 41596 12081 41602
rect 2314 41538 2320 41590
rect 2372 41538 2378 41590
rect 3878 41538 3884 41590
rect 3936 41538 3942 41590
rect 4154 41587 4160 41590
rect 4148 41541 4160 41587
rect 4212 41578 4218 41590
rect 4212 41550 4248 41578
rect 4154 41538 4160 41541
rect 4212 41538 4218 41550
rect 11698 41538 11704 41590
rect 11756 41538 11762 41590
rect 12023 41562 12035 41596
rect 12069 41593 12081 41596
rect 12437 41596 12495 41602
rect 12069 41590 12388 41593
rect 12069 41565 12348 41590
rect 12069 41562 12081 41565
rect 12023 41556 12081 41562
rect 12342 41538 12348 41565
rect 12400 41538 12406 41590
rect 12437 41562 12449 41596
rect 12483 41593 12495 41596
rect 12805 41596 12863 41602
rect 12805 41593 12817 41596
rect 12483 41565 12817 41593
rect 12483 41562 12495 41565
rect 12437 41556 12495 41562
rect 12805 41562 12817 41565
rect 12851 41593 12863 41596
rect 12894 41593 12900 41605
rect 12851 41565 12900 41593
rect 12851 41562 12863 41565
rect 12805 41556 12863 41562
rect 12894 41553 12900 41565
rect 12952 41553 12958 41605
rect 12986 41553 12992 41605
rect 13044 41553 13050 41605
rect 13725 41575 13737 41609
rect 13771 41606 13783 41609
rect 13814 41606 13820 41618
rect 13771 41578 13820 41606
rect 13771 41575 13783 41578
rect 13725 41569 13783 41575
rect 13814 41566 13820 41578
rect 13872 41566 13878 41618
rect 14093 41596 14151 41602
rect 13998 41538 14004 41590
rect 14056 41578 14062 41590
rect 14093 41578 14105 41596
rect 14056 41562 14105 41578
rect 14139 41562 14151 41596
rect 14056 41556 14151 41562
rect 14056 41550 14136 41556
rect 14056 41538 14062 41550
rect 14182 41538 14188 41590
rect 14240 41578 14246 41590
rect 15102 41578 15108 41607
rect 14240 41555 15108 41578
rect 15160 41555 15166 41607
rect 15378 41606 15384 41658
rect 15436 41606 15442 41658
rect 16206 41606 16212 41658
rect 16264 41646 16270 41658
rect 16301 41649 16359 41655
rect 16301 41646 16313 41649
rect 16264 41618 16313 41646
rect 16264 41606 16270 41618
rect 16301 41615 16313 41618
rect 16347 41615 16359 41649
rect 16393 41649 16405 41683
rect 16439 41649 16451 41683
rect 16574 41674 16580 41726
rect 16632 41714 16638 41726
rect 18046 41714 18052 41726
rect 16632 41686 18052 41714
rect 16632 41674 16638 41686
rect 16960 41658 16988 41686
rect 18046 41674 18052 41686
rect 18104 41674 18110 41726
rect 16393 41643 16451 41649
rect 16301 41609 16359 41615
rect 16850 41606 16856 41658
rect 16908 41606 16914 41658
rect 16942 41606 16948 41658
rect 17000 41606 17006 41658
rect 17957 41649 18015 41655
rect 17957 41615 17969 41649
rect 18003 41646 18015 41649
rect 18064 41646 18092 41674
rect 18003 41618 18092 41646
rect 18003 41615 18015 41618
rect 17957 41609 18015 41615
rect 19242 41606 19248 41658
rect 19300 41606 19306 41658
rect 19444 41621 19472 41754
rect 20990 41742 20996 41794
rect 21048 41782 21054 41794
rect 21591 41785 21649 41791
rect 21591 41782 21603 41785
rect 21048 41754 21603 41782
rect 21048 41742 21054 41754
rect 21591 41751 21603 41754
rect 21637 41751 21649 41785
rect 25682 41752 25688 41804
rect 25740 41752 25746 41804
rect 25869 41785 25927 41791
rect 21591 41745 21649 41751
rect 25869 41751 25881 41785
rect 25915 41782 25927 41785
rect 26786 41782 26792 41794
rect 25915 41754 26792 41782
rect 25915 41751 25927 41754
rect 25869 41745 25927 41751
rect 26786 41742 26792 41754
rect 26844 41742 26850 41794
rect 21082 41674 21088 41726
rect 21140 41714 21146 41726
rect 21140 41686 22232 41714
rect 21140 41674 21146 41686
rect 19429 41615 19487 41621
rect 15551 41593 15609 41599
rect 15551 41590 15563 41593
rect 15488 41562 15563 41590
rect 14240 41550 15148 41555
rect 14240 41538 14246 41550
rect 3050 41470 3056 41522
rect 3108 41470 3114 41522
rect 5258 41470 5264 41522
rect 5316 41470 5322 41522
rect 11882 41470 11888 41522
rect 11940 41510 11946 41522
rect 13173 41513 13231 41519
rect 13173 41510 13185 41513
rect 11940 41482 13185 41510
rect 11940 41470 11946 41482
rect 13173 41479 13185 41482
rect 13219 41510 13231 41513
rect 13262 41510 13268 41522
rect 13219 41482 13268 41510
rect 13219 41479 13231 41482
rect 13173 41473 13231 41479
rect 13262 41470 13268 41482
rect 13320 41470 13326 41522
rect 13630 41470 13636 41522
rect 13688 41470 13694 41522
rect 13722 41470 13728 41522
rect 13780 41510 13786 41522
rect 15488 41510 15516 41562
rect 15551 41559 15563 41562
rect 15597 41559 15609 41593
rect 17129 41593 17187 41599
rect 17129 41590 17141 41593
rect 17175 41590 17187 41593
rect 18127 41593 18185 41599
rect 18127 41590 18139 41593
rect 15551 41553 15609 41559
rect 17126 41538 17132 41590
rect 17184 41538 17190 41590
rect 17586 41578 17592 41590
rect 17236 41550 17592 41578
rect 17236 41522 17264 41550
rect 17586 41538 17592 41550
rect 17644 41538 17650 41590
rect 17678 41538 17684 41590
rect 17736 41578 17742 41590
rect 18064 41578 18139 41590
rect 17736 41562 18139 41578
rect 17736 41550 18092 41562
rect 18127 41559 18139 41562
rect 18173 41559 18185 41593
rect 19429 41581 19441 41615
rect 19475 41581 19487 41615
rect 19702 41606 19708 41658
rect 19760 41606 19766 41658
rect 22204 41655 22232 41686
rect 22278 41674 22284 41726
rect 22336 41714 22342 41726
rect 22373 41717 22431 41723
rect 22373 41714 22385 41717
rect 22336 41686 22385 41714
rect 22336 41674 22342 41686
rect 22373 41683 22385 41686
rect 22419 41683 22431 41717
rect 22373 41677 22431 41683
rect 22189 41649 22247 41655
rect 22002 41615 22060 41621
rect 22002 41612 22014 41615
rect 19429 41575 19487 41581
rect 21358 41578 21364 41590
rect 18127 41553 18185 41559
rect 21192 41550 21364 41578
rect 17736 41538 17742 41550
rect 13780 41482 15516 41510
rect 13780 41470 13786 41482
rect 15746 41470 15752 41522
rect 15804 41470 15810 41522
rect 15838 41470 15844 41522
rect 15896 41510 15902 41522
rect 16669 41513 16727 41519
rect 16669 41510 16681 41513
rect 15896 41482 16681 41510
rect 15896 41470 15902 41482
rect 16669 41479 16681 41482
rect 16715 41510 16727 41513
rect 17218 41510 17224 41522
rect 16715 41482 17224 41510
rect 16715 41479 16727 41482
rect 16669 41473 16727 41479
rect 17218 41470 17224 41482
rect 17276 41470 17282 41522
rect 17313 41513 17371 41519
rect 17313 41479 17325 41513
rect 17359 41510 17371 41513
rect 17770 41510 17776 41522
rect 17359 41482 17776 41510
rect 17359 41479 17371 41482
rect 17313 41473 17371 41479
rect 17770 41470 17776 41482
rect 17828 41470 17834 41522
rect 18325 41513 18383 41519
rect 18325 41479 18337 41513
rect 18371 41510 18383 41513
rect 19242 41510 19248 41522
rect 18371 41482 19248 41510
rect 18371 41479 18383 41482
rect 18325 41473 18383 41479
rect 19242 41470 19248 41482
rect 19300 41470 19306 41522
rect 19610 41470 19616 41522
rect 19668 41470 19674 41522
rect 19981 41513 20039 41519
rect 19981 41479 19993 41513
rect 20027 41510 20039 41513
rect 20162 41510 20168 41522
rect 20027 41482 20168 41510
rect 20027 41479 20039 41482
rect 19981 41473 20039 41479
rect 20162 41470 20168 41482
rect 20220 41470 20226 41522
rect 21192 41496 21220 41550
rect 21358 41538 21364 41550
rect 21416 41538 21422 41590
rect 21450 41538 21456 41590
rect 21508 41578 21514 41590
rect 21744 41584 22014 41612
rect 21744 41578 21772 41584
rect 21508 41550 21772 41578
rect 22002 41581 22014 41584
rect 22048 41581 22060 41615
rect 22189 41615 22201 41649
rect 22235 41615 22247 41649
rect 22189 41609 22247 41615
rect 22002 41575 22060 41581
rect 22462 41553 22468 41605
rect 22520 41553 22526 41605
rect 22649 41596 22707 41602
rect 22649 41562 22661 41596
rect 22695 41578 22707 41596
rect 23474 41578 23480 41590
rect 22695 41562 23480 41578
rect 22649 41556 23480 41562
rect 22664 41550 23480 41556
rect 21508 41538 21514 41550
rect 23474 41538 23480 41550
rect 23532 41538 23538 41590
rect 25406 41566 25412 41618
rect 25464 41566 25470 41618
rect 21818 41470 21824 41522
rect 21876 41470 21882 41522
rect 552 41370 31808 41392
rect 552 41318 8172 41370
rect 8224 41318 8236 41370
rect 8288 41318 8300 41370
rect 8352 41318 8364 41370
rect 8416 41318 8428 41370
rect 8480 41318 15946 41370
rect 15998 41318 16010 41370
rect 16062 41318 16074 41370
rect 16126 41318 16138 41370
rect 16190 41318 16202 41370
rect 16254 41318 23720 41370
rect 23772 41318 23784 41370
rect 23836 41318 23848 41370
rect 23900 41318 23912 41370
rect 23964 41318 23976 41370
rect 24028 41318 31494 41370
rect 31546 41318 31558 41370
rect 31610 41318 31622 41370
rect 31674 41318 31686 41370
rect 31738 41318 31750 41370
rect 31802 41318 31808 41370
rect 552 41296 31808 41318
rect 2130 41241 2194 41250
rect 2130 41207 2145 41241
rect 2179 41207 2194 41241
rect 2130 41198 2194 41207
rect 2501 41241 2559 41247
rect 2501 41207 2513 41241
rect 2547 41238 2559 41241
rect 3418 41238 3424 41250
rect 2547 41210 3424 41238
rect 2547 41207 2559 41210
rect 2501 41201 2559 41207
rect 2314 41062 2320 41114
rect 2372 41102 2378 41114
rect 2516 41102 2544 41201
rect 3418 41198 3424 41210
rect 3476 41198 3482 41250
rect 4338 41241 4402 41250
rect 4338 41207 4353 41241
rect 4387 41207 4402 41241
rect 4338 41198 4402 41207
rect 6546 41198 6552 41250
rect 6604 41198 6610 41250
rect 8018 41198 8024 41250
rect 8076 41198 8082 41250
rect 11790 41198 11796 41250
rect 11848 41198 11854 41250
rect 14826 41238 14832 41250
rect 11900 41210 14832 41238
rect 3050 41130 3056 41182
rect 3108 41170 3114 41182
rect 3614 41173 3672 41179
rect 3614 41170 3626 41173
rect 3108 41142 3626 41170
rect 3108 41130 3114 41142
rect 3614 41139 3626 41142
rect 3660 41139 3672 41173
rect 3614 41133 3672 41139
rect 2372 41074 2544 41102
rect 2372 41062 2378 41074
rect 3878 41062 3884 41114
rect 3936 41062 3942 41114
rect 4522 41062 4528 41114
rect 4580 41102 4586 41114
rect 5258 41102 5264 41114
rect 4580 41074 5264 41102
rect 4580 41062 4586 41074
rect 5258 41062 5264 41074
rect 5316 41062 5322 41114
rect 6730 41062 6736 41114
rect 6788 41062 6794 41114
rect 8205 41105 8263 41111
rect 8205 41071 8217 41105
rect 8251 41102 8263 41105
rect 11900 41102 11928 41210
rect 14826 41198 14832 41210
rect 14884 41198 14890 41250
rect 15120 41210 15516 41238
rect 12342 41170 12348 41182
rect 12268 41142 12348 41170
rect 8251 41074 11928 41102
rect 11977 41126 12035 41132
rect 11977 41092 11989 41126
rect 12023 41123 12035 41126
rect 12161 41126 12219 41132
rect 12023 41095 12112 41123
rect 12023 41092 12035 41095
rect 11977 41086 12035 41092
rect 8251 41071 8263 41074
rect 8205 41065 8263 41071
rect 12084 41034 12112 41095
rect 12161 41092 12173 41126
rect 12207 41123 12219 41126
rect 12268 41123 12296 41142
rect 12342 41130 12348 41142
rect 12400 41170 12406 41182
rect 12400 41142 12756 41170
rect 12400 41130 12406 41142
rect 12207 41095 12296 41123
rect 12728 41123 12756 41142
rect 12805 41126 12863 41132
rect 12805 41123 12817 41126
rect 12207 41092 12219 41095
rect 12161 41086 12219 41092
rect 12526 41062 12532 41114
rect 12584 41062 12590 41114
rect 12618 41062 12624 41114
rect 12676 41111 12682 41114
rect 12676 41105 12696 41111
rect 12684 41071 12696 41105
rect 12728 41095 12817 41123
rect 12805 41092 12817 41095
rect 12851 41092 12863 41126
rect 12805 41086 12863 41092
rect 12676 41065 12696 41071
rect 12912 41074 13584 41102
rect 13630 41082 13636 41134
rect 13688 41082 13694 41134
rect 13814 41130 13820 41182
rect 13872 41170 13878 41182
rect 13872 41145 14135 41170
rect 13872 41142 14150 41145
rect 13872 41130 13878 41142
rect 14092 41139 14150 41142
rect 14092 41105 14104 41139
rect 14138 41105 14150 41139
rect 14274 41130 14280 41182
rect 14332 41130 14338 41182
rect 14092 41099 14150 41105
rect 12676 41062 12682 41065
rect 12912 41034 12940 41074
rect 12084 41006 12940 41034
rect 13556 41034 13584 41074
rect 14366 41062 14372 41114
rect 14424 41062 14430 41114
rect 14550 41083 14556 41135
rect 14608 41123 14614 41135
rect 15120 41132 15148 41210
rect 15488 41170 15516 41210
rect 15562 41198 15568 41250
rect 15620 41238 15626 41250
rect 15657 41241 15715 41247
rect 15657 41238 15669 41241
rect 15620 41210 15669 41238
rect 15620 41198 15626 41210
rect 15657 41207 15669 41210
rect 15703 41207 15715 41241
rect 16666 41238 16672 41250
rect 15657 41201 15715 41207
rect 16408 41210 16672 41238
rect 15838 41170 15844 41182
rect 15488 41142 15844 41170
rect 15105 41126 15163 41132
rect 14608 41095 15056 41123
rect 14608 41083 14614 41095
rect 13817 41037 13875 41043
rect 13817 41034 13829 41037
rect 13556 41006 13829 41034
rect 13817 41003 13829 41006
rect 13863 41034 13875 41037
rect 13906 41034 13912 41046
rect 13863 41006 13912 41034
rect 13863 41003 13875 41006
rect 13817 40997 13875 41003
rect 13906 40994 13912 41006
rect 13964 40994 13970 41046
rect 15028 41034 15056 41095
rect 15105 41092 15117 41126
rect 15151 41092 15163 41126
rect 15335 41126 15393 41132
rect 15838 41130 15844 41142
rect 15896 41130 15902 41182
rect 16408 41132 16436 41210
rect 16666 41198 16672 41210
rect 16724 41198 16730 41250
rect 17052 41210 17908 41238
rect 15335 41123 15347 41126
rect 15105 41086 15163 41092
rect 15212 41095 15347 41123
rect 15212 41046 15240 41095
rect 15335 41092 15347 41095
rect 15381 41092 15393 41126
rect 15933 41126 15991 41132
rect 15335 41086 15393 41092
rect 15470 41062 15476 41114
rect 15528 41102 15534 41114
rect 15528 41074 15884 41102
rect 15933 41092 15945 41126
rect 15979 41123 15991 41126
rect 16393 41126 16451 41132
rect 16393 41123 16405 41126
rect 15979 41095 16405 41123
rect 15979 41092 15991 41095
rect 15933 41086 15991 41092
rect 16393 41092 16405 41095
rect 16439 41092 16451 41126
rect 16393 41086 16451 41092
rect 16482 41083 16488 41135
rect 16540 41123 16546 41135
rect 16577 41126 16635 41132
rect 16577 41123 16589 41126
rect 16540 41095 16589 41123
rect 16540 41083 16546 41095
rect 16577 41092 16589 41095
rect 16623 41123 16635 41126
rect 16945 41126 17003 41132
rect 16945 41123 16957 41126
rect 16623 41095 16957 41123
rect 16623 41092 16635 41095
rect 16577 41086 16635 41092
rect 16945 41092 16957 41095
rect 16991 41092 17003 41126
rect 16945 41086 17003 41092
rect 15528 41062 15534 41074
rect 15194 41034 15200 41046
rect 15028 41006 15200 41034
rect 15194 40994 15200 41006
rect 15252 40994 15258 41046
rect 15856 40966 15884 41074
rect 16114 40994 16120 41046
rect 16172 40994 16178 41046
rect 17052 41034 17080 41210
rect 17218 41083 17224 41135
rect 17276 41123 17282 41135
rect 17359 41126 17417 41132
rect 17494 41130 17500 41182
rect 17552 41170 17558 41182
rect 17681 41173 17739 41179
rect 17681 41170 17693 41173
rect 17552 41142 17693 41170
rect 17552 41130 17558 41142
rect 17681 41139 17693 41142
rect 17727 41139 17739 41173
rect 17681 41133 17739 41139
rect 17359 41123 17371 41126
rect 17276 41095 17371 41123
rect 17276 41083 17282 41095
rect 17359 41092 17371 41095
rect 17405 41092 17417 41126
rect 17359 41086 17417 41092
rect 17770 41062 17776 41114
rect 17828 41062 17834 41114
rect 17880 41102 17908 41210
rect 17954 41198 17960 41250
rect 18012 41198 18018 41250
rect 20441 41241 20499 41247
rect 20441 41207 20453 41241
rect 20487 41238 20499 41241
rect 20622 41238 20628 41250
rect 20487 41210 20628 41238
rect 20487 41207 20499 41210
rect 20441 41201 20499 41207
rect 20622 41198 20628 41210
rect 20680 41198 20686 41250
rect 22189 41241 22247 41247
rect 20824 41210 22140 41238
rect 19242 41130 19248 41182
rect 19300 41130 19306 41182
rect 19352 41142 20668 41170
rect 19352 41102 19380 41142
rect 17880 41074 19380 41102
rect 19610 41062 19616 41114
rect 19668 41102 19674 41114
rect 20257 41105 20315 41111
rect 20257 41102 20269 41105
rect 19668 41074 20269 41102
rect 19668 41062 19674 41074
rect 20257 41071 20269 41074
rect 20303 41071 20315 41105
rect 20640 41102 20668 41142
rect 20714 41130 20720 41182
rect 20772 41130 20778 41182
rect 20824 41102 20852 41210
rect 21818 41130 21824 41182
rect 21876 41130 21882 41182
rect 20640 41074 20852 41102
rect 20257 41065 20315 41071
rect 20898 41062 20904 41114
rect 20956 41102 20962 41114
rect 22005 41105 22063 41111
rect 22005 41102 22017 41105
rect 20956 41074 22017 41102
rect 20956 41062 20962 41074
rect 22005 41071 22017 41074
rect 22051 41071 22063 41105
rect 22112 41102 22140 41210
rect 22189 41207 22201 41241
rect 22235 41207 22247 41241
rect 22189 41201 22247 41207
rect 22204 41170 22232 41201
rect 22830 41170 22836 41182
rect 22204 41142 22836 41170
rect 22830 41130 22836 41142
rect 22888 41130 22894 41182
rect 23469 41129 23527 41135
rect 30190 41130 30196 41182
rect 30248 41130 30254 41182
rect 23469 41126 23481 41129
rect 23216 41102 23481 41126
rect 22112 41098 23481 41102
rect 22112 41074 23244 41098
rect 23469 41095 23481 41098
rect 23515 41095 23527 41129
rect 30480 41122 30538 41128
rect 23469 41089 23527 41095
rect 22005 41065 22063 41071
rect 23566 41062 23572 41114
rect 23624 41062 23630 41114
rect 30480 41088 30492 41122
rect 30526 41119 30538 41122
rect 30742 41119 30748 41131
rect 30526 41091 30748 41119
rect 30526 41088 30538 41091
rect 30480 41082 30538 41088
rect 30742 41079 30748 41091
rect 30800 41079 30806 41131
rect 16960 41006 17080 41034
rect 20993 41037 21051 41043
rect 16960 40966 16988 41006
rect 20993 41003 21005 41037
rect 21039 41034 21051 41037
rect 22094 41034 22100 41046
rect 21039 41006 22100 41034
rect 21039 41003 21051 41006
rect 20993 40997 21051 41003
rect 22094 40994 22100 41006
rect 22152 40994 22158 41046
rect 27246 41034 27252 41046
rect 22204 41006 27252 41034
rect 15856 40938 16988 40966
rect 19518 40926 19524 40978
rect 19576 40926 19582 40978
rect 21729 40969 21787 40975
rect 21729 40935 21741 40969
rect 21775 40966 21787 40969
rect 22204 40966 22232 41006
rect 27246 40994 27252 41006
rect 27304 40994 27310 41046
rect 21775 40938 22232 40966
rect 21775 40935 21787 40938
rect 21729 40929 21787 40935
rect 22278 40926 22284 40978
rect 22336 40966 22342 40978
rect 25774 40966 25780 40978
rect 22336 40938 25780 40966
rect 22336 40926 22342 40938
rect 25774 40926 25780 40938
rect 25832 40926 25838 40978
rect 200 40826 31648 40848
rect 200 40774 206 40826
rect 514 40774 4285 40826
rect 4337 40774 4349 40826
rect 4401 40774 4413 40826
rect 4465 40774 4477 40826
rect 4529 40774 4541 40826
rect 4593 40774 12059 40826
rect 12111 40774 12123 40826
rect 12175 40774 12187 40826
rect 12239 40774 12251 40826
rect 12303 40774 12315 40826
rect 12367 40774 19833 40826
rect 19885 40774 19897 40826
rect 19949 40774 19961 40826
rect 20013 40774 20025 40826
rect 20077 40774 20089 40826
rect 20141 40774 27607 40826
rect 27659 40774 27671 40826
rect 27723 40774 27735 40826
rect 27787 40774 27799 40826
rect 27851 40774 27863 40826
rect 27915 40774 31648 40826
rect 200 40752 31648 40774
rect 19518 40654 19524 40706
rect 19576 40694 19582 40706
rect 28718 40694 28724 40706
rect 19576 40666 28724 40694
rect 19576 40654 19582 40666
rect 28718 40654 28724 40666
rect 28776 40654 28782 40706
rect 15378 40626 15384 40638
rect 13096 40598 15384 40626
rect 13096 40567 13124 40598
rect 15378 40586 15384 40598
rect 15436 40626 15442 40638
rect 16942 40626 16948 40638
rect 15436 40598 16948 40626
rect 15436 40586 15442 40598
rect 16942 40586 16948 40598
rect 17000 40586 17006 40638
rect 13081 40561 13139 40567
rect 13081 40527 13093 40561
rect 13127 40527 13139 40561
rect 13081 40521 13139 40527
rect 12877 40505 12935 40511
rect 12877 40502 12889 40505
rect 12434 40450 12440 40502
rect 12492 40490 12498 40502
rect 12636 40490 12889 40502
rect 12492 40474 12889 40490
rect 12492 40462 12664 40474
rect 12877 40471 12889 40474
rect 12923 40471 12935 40505
rect 12877 40465 12935 40471
rect 15013 40493 15071 40499
rect 12492 40450 12498 40462
rect 15013 40459 15025 40493
rect 15059 40459 15071 40493
rect 15194 40465 15200 40517
rect 15252 40465 15258 40517
rect 15654 40465 15660 40517
rect 15712 40465 15718 40517
rect 15013 40453 15071 40459
rect 6730 40382 6736 40434
rect 6788 40422 6794 40434
rect 12713 40425 12771 40431
rect 12713 40422 12725 40425
rect 6788 40394 12725 40422
rect 6788 40382 6794 40394
rect 12713 40391 12725 40394
rect 12759 40391 12771 40425
rect 12713 40385 12771 40391
rect 12802 40382 12808 40434
rect 12860 40422 12866 40434
rect 15028 40422 15056 40453
rect 15746 40450 15752 40502
rect 15804 40490 15810 40502
rect 16117 40493 16175 40499
rect 16117 40490 16129 40493
rect 15804 40462 16129 40490
rect 15804 40450 15810 40462
rect 16117 40459 16129 40462
rect 16163 40459 16175 40493
rect 16117 40453 16175 40459
rect 12860 40394 15056 40422
rect 16301 40425 16359 40431
rect 12860 40382 12866 40394
rect 16301 40391 16313 40425
rect 16347 40422 16359 40425
rect 16942 40422 16948 40434
rect 16347 40394 16948 40422
rect 16347 40391 16359 40394
rect 16301 40385 16359 40391
rect 16942 40382 16948 40394
rect 17000 40382 17006 40434
rect 552 40282 31808 40304
rect 552 40230 8172 40282
rect 8224 40230 8236 40282
rect 8288 40230 8300 40282
rect 8352 40230 8364 40282
rect 8416 40230 8428 40282
rect 8480 40230 15946 40282
rect 15998 40230 16010 40282
rect 16062 40230 16074 40282
rect 16126 40230 16138 40282
rect 16190 40230 16202 40282
rect 16254 40230 23720 40282
rect 23772 40230 23784 40282
rect 23836 40230 23848 40282
rect 23900 40230 23912 40282
rect 23964 40230 23976 40282
rect 24028 40230 31494 40282
rect 31546 40230 31558 40282
rect 31610 40230 31622 40282
rect 31674 40230 31686 40282
rect 31738 40230 31750 40282
rect 31802 40230 31808 40282
rect 552 40208 31808 40230
rect 8128 40048 10522 40056
rect 8128 39968 8148 40048
rect 8502 40040 10522 40048
rect 10502 39976 10522 40040
rect 8502 39968 10522 39976
rect 8128 39960 10522 39968
rect 9630 39800 9714 39960
rect 1051 39792 1157 39799
rect 1051 39740 1058 39792
rect 1150 39740 1157 39792
rect 1051 39733 1157 39740
rect 9134 39728 10214 39800
rect 18202 39790 18310 39800
rect 18202 39738 18212 39790
rect 18300 39738 18310 39790
rect 18202 39728 18310 39738
rect 31498 39758 31792 39764
rect 9630 39560 9714 39728
rect 31498 39560 31518 39758
rect 220 39553 31518 39560
rect 220 39489 239 39553
rect 220 39488 31518 39489
rect 31772 39488 31792 39758
rect 220 39482 31792 39488
<< via1 >>
rect 15752 44734 15804 44786
rect 23296 44734 23348 44786
rect 23480 44734 23532 44786
rect 30380 44734 30432 44786
rect 8172 44582 8224 44634
rect 8236 44582 8288 44634
rect 8300 44582 8352 44634
rect 8364 44582 8416 44634
rect 8428 44582 8480 44634
rect 15946 44582 15998 44634
rect 16010 44582 16062 44634
rect 16074 44582 16126 44634
rect 16138 44582 16190 44634
rect 16202 44582 16254 44634
rect 23720 44582 23772 44634
rect 23784 44582 23836 44634
rect 23848 44582 23900 44634
rect 23912 44582 23964 44634
rect 23976 44582 24028 44634
rect 31494 44582 31546 44634
rect 31558 44582 31610 44634
rect 31622 44582 31674 44634
rect 31686 44582 31738 44634
rect 31750 44582 31802 44634
rect 848 44505 900 44514
rect 848 44471 857 44505
rect 857 44471 891 44505
rect 891 44471 900 44505
rect 848 44462 900 44471
rect 1584 44505 1636 44514
rect 1584 44471 1593 44505
rect 1593 44471 1627 44505
rect 1627 44471 1636 44505
rect 1584 44462 1636 44471
rect 2320 44505 2372 44514
rect 2320 44471 2329 44505
rect 2329 44471 2363 44505
rect 2363 44471 2372 44505
rect 2320 44462 2372 44471
rect 3240 44505 3292 44514
rect 3240 44471 3249 44505
rect 3249 44471 3283 44505
rect 3283 44471 3292 44505
rect 3240 44462 3292 44471
rect 3792 44505 3844 44514
rect 3792 44471 3801 44505
rect 3801 44471 3835 44505
rect 3835 44471 3844 44505
rect 3792 44462 3844 44471
rect 4528 44505 4580 44514
rect 4528 44471 4537 44505
rect 4537 44471 4571 44505
rect 4571 44471 4580 44505
rect 4528 44462 4580 44471
rect 5264 44505 5316 44514
rect 5264 44471 5273 44505
rect 5273 44471 5307 44505
rect 5307 44471 5316 44505
rect 5264 44462 5316 44471
rect 6000 44505 6052 44514
rect 6000 44471 6009 44505
rect 6009 44471 6043 44505
rect 6043 44471 6052 44505
rect 6000 44462 6052 44471
rect 9680 44394 9732 44446
rect 13912 44462 13964 44514
rect 12624 44347 12676 44399
rect 13360 44394 13412 44446
rect 14096 44505 14148 44514
rect 14096 44471 14105 44505
rect 14105 44471 14139 44505
rect 14139 44471 14148 44505
rect 14096 44462 14148 44471
rect 15660 44462 15712 44514
rect 14372 44394 14424 44446
rect 13544 44326 13596 44378
rect 12532 44233 12584 44242
rect 12532 44199 12541 44233
rect 12541 44199 12575 44233
rect 12575 44199 12584 44233
rect 12532 44190 12584 44199
rect 13268 44258 13320 44310
rect 13360 44258 13412 44310
rect 13820 44385 13872 44394
rect 13820 44351 13829 44385
rect 13829 44351 13863 44385
rect 13863 44351 13872 44385
rect 13820 44342 13872 44351
rect 14280 44369 14332 44378
rect 14280 44335 14289 44369
rect 14289 44335 14323 44369
rect 14323 44335 14332 44369
rect 14280 44326 14332 44335
rect 15568 44350 15620 44402
rect 15752 44403 15804 44412
rect 15752 44369 15761 44403
rect 15761 44369 15795 44403
rect 15795 44369 15804 44403
rect 15752 44360 15804 44369
rect 16304 44347 16356 44399
rect 17868 44462 17920 44514
rect 19156 44462 19208 44514
rect 16856 44390 16908 44399
rect 16856 44356 16865 44390
rect 16865 44356 16899 44390
rect 16899 44356 16908 44390
rect 16856 44347 16908 44356
rect 17040 44437 17092 44446
rect 17040 44403 17049 44437
rect 17049 44403 17083 44437
rect 17083 44403 17092 44437
rect 17040 44394 17092 44403
rect 19616 44462 19668 44514
rect 17224 44326 17276 44378
rect 21824 44394 21876 44446
rect 18972 44326 19024 44378
rect 19064 44334 19116 44386
rect 19248 44377 19300 44386
rect 19248 44343 19257 44377
rect 19257 44343 19291 44377
rect 19291 44343 19300 44377
rect 19248 44334 19300 44343
rect 21916 44369 21968 44378
rect 21916 44335 21925 44369
rect 21925 44335 21959 44369
rect 21959 44335 21968 44369
rect 21916 44326 21968 44335
rect 14924 44258 14976 44310
rect 15476 44258 15528 44310
rect 21732 44258 21784 44310
rect 22100 44326 22152 44378
rect 23020 44326 23072 44378
rect 26516 44394 26568 44446
rect 31116 44462 31168 44514
rect 23204 44369 23256 44378
rect 23204 44335 23213 44369
rect 23213 44335 23247 44369
rect 23247 44335 23256 44369
rect 23204 44326 23256 44335
rect 24124 44258 24176 44310
rect 25228 44369 25280 44378
rect 25228 44335 25237 44369
rect 25237 44335 25271 44369
rect 25271 44335 25280 44369
rect 25228 44326 25280 44335
rect 25504 44369 25556 44378
rect 25504 44335 25513 44369
rect 25513 44335 25547 44369
rect 25547 44335 25556 44369
rect 25504 44326 25556 44335
rect 26792 44369 26844 44378
rect 26792 44335 26801 44369
rect 26801 44335 26835 44369
rect 26835 44335 26844 44369
rect 26792 44326 26844 44335
rect 27988 44326 28040 44378
rect 28632 44369 28684 44378
rect 28632 44335 28641 44369
rect 28641 44335 28675 44369
rect 28675 44335 28684 44369
rect 28632 44326 28684 44335
rect 13176 44190 13228 44242
rect 13820 44233 13872 44242
rect 13820 44199 13829 44233
rect 13829 44199 13863 44233
rect 13863 44199 13872 44233
rect 13820 44190 13872 44199
rect 16396 44190 16448 44242
rect 16580 44190 16632 44242
rect 19340 44233 19392 44242
rect 19340 44199 19349 44233
rect 19349 44199 19383 44233
rect 19383 44199 19392 44233
rect 19340 44190 19392 44199
rect 21640 44190 21692 44242
rect 22008 44190 22060 44242
rect 22100 44233 22152 44242
rect 22100 44199 22109 44233
rect 22109 44199 22143 44233
rect 22143 44199 22152 44233
rect 22100 44190 22152 44199
rect 26240 44258 26292 44310
rect 27528 44258 27580 44310
rect 29184 44258 29236 44310
rect 30472 44326 30524 44378
rect 30564 44326 30616 44378
rect 30840 44258 30892 44310
rect 26608 44233 26660 44242
rect 26608 44199 26617 44233
rect 26617 44199 26651 44233
rect 26651 44199 26660 44233
rect 26608 44190 26660 44199
rect 27068 44190 27120 44242
rect 29460 44190 29512 44242
rect 30564 44233 30616 44242
rect 30564 44199 30573 44233
rect 30573 44199 30607 44233
rect 30607 44199 30616 44233
rect 30564 44190 30616 44199
rect 206 44038 514 44090
rect 4285 44038 4337 44090
rect 4349 44038 4401 44090
rect 4413 44038 4465 44090
rect 4477 44038 4529 44090
rect 4541 44038 4593 44090
rect 12059 44038 12111 44090
rect 12123 44038 12175 44090
rect 12187 44038 12239 44090
rect 12251 44038 12303 44090
rect 12315 44038 12367 44090
rect 19833 44038 19885 44090
rect 19897 44038 19949 44090
rect 19961 44038 20013 44090
rect 20025 44038 20077 44090
rect 20089 44038 20141 44090
rect 27607 44038 27659 44090
rect 27671 44038 27723 44090
rect 27735 44038 27787 44090
rect 27799 44038 27851 44090
rect 27863 44038 27915 44090
rect 11336 43714 11388 43766
rect 11520 43757 11572 43766
rect 11520 43723 11529 43757
rect 11529 43723 11563 43757
rect 11563 43723 11572 43757
rect 11520 43714 11572 43723
rect 17224 43961 17276 43970
rect 17224 43927 17233 43961
rect 17233 43927 17267 43961
rect 17267 43927 17276 43961
rect 17224 43918 17276 43927
rect 22008 43918 22060 43970
rect 23664 43961 23716 43970
rect 23664 43927 23673 43961
rect 23673 43927 23707 43961
rect 23707 43927 23716 43961
rect 23664 43918 23716 43927
rect 27528 43918 27580 43970
rect 11244 43689 11296 43698
rect 11244 43655 11253 43689
rect 11253 43655 11287 43689
rect 11287 43655 11296 43689
rect 11244 43646 11296 43655
rect 14004 43782 14056 43834
rect 14188 43714 14240 43766
rect 14372 43772 14424 43781
rect 14372 43738 14381 43772
rect 14381 43738 14415 43772
rect 14415 43738 14424 43772
rect 14372 43729 14424 43738
rect 13176 43646 13228 43698
rect 14004 43646 14056 43698
rect 14464 43646 14516 43698
rect 14740 43689 14792 43698
rect 14740 43655 14749 43689
rect 14749 43655 14783 43689
rect 14783 43655 14792 43689
rect 14740 43646 14792 43655
rect 15384 43714 15436 43766
rect 15476 43757 15528 43766
rect 15476 43723 15485 43757
rect 15485 43723 15519 43757
rect 15519 43723 15528 43757
rect 15476 43714 15528 43723
rect 15568 43714 15620 43766
rect 15200 43646 15252 43698
rect 15292 43646 15344 43698
rect 16580 43714 16632 43766
rect 19064 43850 19116 43902
rect 19892 43850 19944 43902
rect 21916 43850 21968 43902
rect 23204 43850 23256 43902
rect 28080 43918 28132 43970
rect 28908 43918 28960 43970
rect 30380 43961 30432 43970
rect 30380 43927 30389 43961
rect 30389 43927 30423 43961
rect 30423 43927 30432 43961
rect 30380 43918 30432 43927
rect 30472 43918 30524 43970
rect 17408 43825 17460 43834
rect 17408 43791 17417 43825
rect 17417 43791 17451 43825
rect 17451 43791 17460 43825
rect 17408 43782 17460 43791
rect 17960 43782 18012 43834
rect 19708 43782 19760 43834
rect 17592 43772 17644 43781
rect 17592 43738 17601 43772
rect 17601 43738 17635 43772
rect 17635 43738 17644 43772
rect 17592 43729 17644 43738
rect 17868 43772 17920 43781
rect 17868 43738 17877 43772
rect 17877 43738 17911 43772
rect 17911 43738 17920 43772
rect 17868 43729 17920 43738
rect 18788 43646 18840 43698
rect 19616 43757 19668 43766
rect 19616 43723 19625 43757
rect 19625 43723 19659 43757
rect 19659 43723 19668 43757
rect 19616 43714 19668 43723
rect 19892 43757 19944 43766
rect 19892 43723 19901 43757
rect 19901 43723 19935 43757
rect 19935 43723 19944 43757
rect 19892 43714 19944 43723
rect 21640 43782 21692 43834
rect 22928 43825 22980 43834
rect 22928 43791 22937 43825
rect 22937 43791 22971 43825
rect 22971 43791 22980 43825
rect 22928 43782 22980 43791
rect 22652 43757 22704 43766
rect 22652 43723 22670 43757
rect 22670 43723 22704 43757
rect 22652 43714 22704 43723
rect 23388 43757 23440 43766
rect 23388 43723 23397 43757
rect 23397 43723 23431 43757
rect 23431 43723 23440 43757
rect 23388 43714 23440 43723
rect 31116 43825 31168 43834
rect 31116 43791 31125 43825
rect 31125 43791 31159 43825
rect 31159 43791 31168 43825
rect 31116 43782 31168 43791
rect 24584 43757 24636 43766
rect 24584 43723 24596 43757
rect 24596 43723 24636 43757
rect 22928 43646 22980 43698
rect 23020 43689 23072 43698
rect 23020 43655 23029 43689
rect 23029 43655 23063 43689
rect 23063 43655 23072 43689
rect 23020 43646 23072 43655
rect 23204 43646 23256 43698
rect 23572 43646 23624 43698
rect 24584 43714 24636 43723
rect 24400 43646 24452 43698
rect 26884 43757 26936 43766
rect 26884 43723 26918 43757
rect 26918 43723 26936 43757
rect 25504 43646 25556 43698
rect 26884 43714 26936 43723
rect 29000 43757 29052 43766
rect 29000 43723 29009 43757
rect 29009 43723 29043 43757
rect 29043 43723 29052 43757
rect 29000 43714 29052 43723
rect 29276 43757 29328 43766
rect 29276 43723 29310 43757
rect 29310 43723 29328 43757
rect 29276 43714 29328 43723
rect 27988 43689 28040 43698
rect 27988 43655 27997 43689
rect 27997 43655 28031 43689
rect 28031 43655 28040 43689
rect 27988 43646 28040 43655
rect 28356 43689 28408 43698
rect 28356 43655 28365 43689
rect 28365 43655 28399 43689
rect 28399 43655 28408 43689
rect 28356 43646 28408 43655
rect 28632 43646 28684 43698
rect 29368 43646 29420 43698
rect 8172 43494 8224 43546
rect 8236 43494 8288 43546
rect 8300 43494 8352 43546
rect 8364 43494 8416 43546
rect 8428 43494 8480 43546
rect 15946 43494 15998 43546
rect 16010 43494 16062 43546
rect 16074 43494 16126 43546
rect 16138 43494 16190 43546
rect 16202 43494 16254 43546
rect 23720 43494 23772 43546
rect 23784 43494 23836 43546
rect 23848 43494 23900 43546
rect 23912 43494 23964 43546
rect 23976 43494 24028 43546
rect 31494 43494 31546 43546
rect 31558 43494 31610 43546
rect 31622 43494 31674 43546
rect 31686 43494 31738 43546
rect 31750 43494 31802 43546
rect 14188 43417 14240 43426
rect 14188 43383 14197 43417
rect 14197 43383 14231 43417
rect 14231 43383 14240 43417
rect 14188 43374 14240 43383
rect 13176 43349 13228 43358
rect 13176 43315 13185 43349
rect 13185 43315 13219 43349
rect 13219 43315 13228 43349
rect 13176 43306 13228 43315
rect 13084 43281 13136 43290
rect 13084 43247 13093 43281
rect 13093 43247 13127 43281
rect 13127 43247 13136 43281
rect 13084 43238 13136 43247
rect 13268 43238 13320 43290
rect 14372 43281 14424 43290
rect 14372 43247 14390 43281
rect 14390 43247 14424 43281
rect 14372 43238 14424 43247
rect 14924 43238 14976 43290
rect 19248 43374 19300 43426
rect 19340 43374 19392 43426
rect 16396 43349 16448 43358
rect 16396 43315 16430 43349
rect 16430 43315 16448 43349
rect 16396 43306 16448 43315
rect 18788 43349 18840 43358
rect 18788 43315 18806 43349
rect 18806 43315 18840 43349
rect 19616 43383 19668 43392
rect 19616 43349 19625 43383
rect 19625 43349 19659 43383
rect 19659 43349 19668 43383
rect 19616 43340 19668 43349
rect 22652 43374 22704 43426
rect 22928 43417 22980 43426
rect 22928 43383 22937 43417
rect 22937 43383 22971 43417
rect 22971 43383 22980 43417
rect 22928 43374 22980 43383
rect 23388 43374 23440 43426
rect 18788 43306 18840 43315
rect 15384 43238 15436 43290
rect 23204 43306 23256 43358
rect 23940 43306 23992 43358
rect 19248 43238 19300 43290
rect 21456 43281 21508 43290
rect 21456 43247 21465 43281
rect 21465 43247 21499 43281
rect 21499 43247 21508 43281
rect 21456 43238 21508 43247
rect 23572 43281 23624 43290
rect 23572 43247 23581 43281
rect 23581 43247 23615 43281
rect 23615 43247 23624 43281
rect 23572 43238 23624 43247
rect 24676 43306 24728 43358
rect 25504 43349 25556 43358
rect 25504 43315 25513 43349
rect 25513 43315 25547 43349
rect 25547 43315 25556 43349
rect 25504 43306 25556 43315
rect 26608 43374 26660 43426
rect 26884 43417 26936 43426
rect 26884 43383 26893 43417
rect 26893 43383 26927 43417
rect 26927 43383 26936 43417
rect 26884 43374 26936 43383
rect 28356 43374 28408 43426
rect 27988 43306 28040 43358
rect 29552 43374 29604 43426
rect 30472 43306 30524 43358
rect 11336 43213 11388 43222
rect 11336 43179 11345 43213
rect 11345 43179 11379 43213
rect 11379 43179 11388 43213
rect 11336 43170 11388 43179
rect 12624 43170 12676 43222
rect 13544 43170 13596 43222
rect 15292 43170 15344 43222
rect 17316 43170 17368 43222
rect 17960 43170 18012 43222
rect 25228 43289 25280 43298
rect 25228 43255 25237 43289
rect 25237 43255 25271 43289
rect 25271 43255 25280 43289
rect 25228 43246 25280 43255
rect 11796 43102 11848 43154
rect 15200 43145 15252 43154
rect 15200 43111 15209 43145
rect 15209 43111 15243 43145
rect 15243 43111 15252 43145
rect 15200 43102 15252 43111
rect 16120 43102 16172 43154
rect 17040 43102 17092 43154
rect 22560 43102 22612 43154
rect 25044 43170 25096 43222
rect 26056 43213 26108 43222
rect 26056 43179 26065 43213
rect 26065 43179 26099 43213
rect 26099 43179 26108 43213
rect 26056 43170 26108 43179
rect 26240 43213 26292 43222
rect 26240 43179 26249 43213
rect 26249 43179 26283 43213
rect 26283 43179 26292 43213
rect 26240 43170 26292 43179
rect 26516 43238 26568 43290
rect 27068 43281 27120 43290
rect 27068 43247 27077 43281
rect 27077 43247 27111 43281
rect 27111 43247 27120 43281
rect 27068 43238 27120 43247
rect 27436 43213 27488 43222
rect 27436 43179 27445 43213
rect 27445 43179 27479 43213
rect 27479 43179 27488 43213
rect 27436 43170 27488 43179
rect 28908 43238 28960 43290
rect 29368 43281 29420 43290
rect 29368 43247 29377 43281
rect 29377 43247 29411 43281
rect 29411 43247 29420 43281
rect 29368 43238 29420 43247
rect 30840 43374 30892 43426
rect 29000 43170 29052 43222
rect 26424 43145 26476 43154
rect 26424 43111 26433 43145
rect 26433 43111 26467 43145
rect 26467 43111 26476 43145
rect 26424 43102 26476 43111
rect 31116 43102 31168 43154
rect 206 42950 514 43002
rect 4285 42950 4337 43002
rect 4349 42950 4401 43002
rect 4413 42950 4465 43002
rect 4477 42950 4529 43002
rect 4541 42950 4593 43002
rect 12059 42950 12111 43002
rect 12123 42950 12175 43002
rect 12187 42950 12239 43002
rect 12251 42950 12303 43002
rect 12315 42950 12367 43002
rect 19833 42950 19885 43002
rect 19897 42950 19949 43002
rect 19961 42950 20013 43002
rect 20025 42950 20077 43002
rect 20089 42950 20141 43002
rect 27607 42950 27659 43002
rect 27671 42950 27723 43002
rect 27735 42950 27787 43002
rect 27799 42950 27851 43002
rect 27863 42950 27915 43002
rect 11152 42873 11204 42882
rect 11152 42839 11161 42873
rect 11161 42839 11195 42873
rect 11195 42839 11204 42873
rect 11152 42830 11204 42839
rect 12440 42830 12492 42882
rect 13084 42830 13136 42882
rect 21456 42830 21508 42882
rect 21824 42830 21876 42882
rect 12624 42762 12676 42814
rect 13360 42762 13412 42814
rect 14924 42694 14976 42746
rect 15016 42694 15068 42746
rect 15384 42762 15436 42814
rect 12532 42626 12584 42678
rect 12164 42601 12216 42610
rect 12164 42567 12173 42601
rect 12173 42567 12207 42601
rect 12207 42567 12216 42601
rect 12164 42558 12216 42567
rect 12348 42558 12400 42610
rect 12992 42669 13044 42678
rect 12992 42635 13001 42669
rect 13001 42635 13035 42669
rect 13035 42635 13044 42669
rect 12992 42626 13044 42635
rect 13084 42626 13136 42678
rect 13452 42641 13504 42693
rect 16948 42694 17000 42746
rect 15200 42626 15252 42678
rect 15292 42669 15344 42678
rect 15292 42635 15301 42669
rect 15301 42635 15335 42669
rect 15335 42635 15344 42669
rect 15292 42626 15344 42635
rect 13544 42558 13596 42610
rect 14188 42601 14240 42610
rect 14188 42567 14197 42601
rect 14197 42567 14231 42601
rect 14231 42567 14240 42601
rect 14188 42558 14240 42567
rect 15384 42558 15436 42610
rect 15660 42626 15712 42678
rect 16304 42684 16356 42693
rect 16304 42650 16313 42684
rect 16313 42650 16347 42684
rect 16347 42650 16356 42684
rect 16304 42641 16356 42650
rect 17316 42558 17368 42610
rect 18236 42601 18288 42610
rect 18236 42567 18245 42601
rect 18245 42567 18279 42601
rect 18279 42567 18288 42601
rect 18236 42558 18288 42567
rect 19616 42694 19668 42746
rect 20904 42694 20956 42746
rect 21088 42694 21140 42746
rect 21824 42737 21876 42746
rect 21824 42703 21833 42737
rect 21833 42703 21867 42737
rect 21867 42703 21876 42737
rect 21824 42694 21876 42703
rect 22560 42737 22612 42746
rect 22560 42703 22569 42737
rect 22569 42703 22603 42737
rect 22603 42703 22612 42737
rect 22560 42694 22612 42703
rect 23480 42694 23532 42746
rect 24124 42762 24176 42814
rect 22376 42626 22428 42678
rect 19892 42558 19944 42610
rect 20812 42601 20864 42610
rect 20812 42567 20821 42601
rect 20821 42567 20855 42601
rect 20855 42567 20864 42601
rect 20812 42558 20864 42567
rect 21180 42558 21232 42610
rect 21456 42558 21508 42610
rect 22744 42601 22796 42610
rect 22744 42567 22753 42601
rect 22753 42567 22787 42601
rect 22787 42567 22796 42601
rect 22744 42558 22796 42567
rect 23020 42558 23072 42610
rect 23204 42669 23256 42678
rect 23204 42635 23213 42669
rect 23213 42635 23247 42669
rect 23247 42635 23256 42669
rect 23204 42626 23256 42635
rect 23480 42601 23532 42610
rect 23480 42567 23489 42601
rect 23489 42567 23523 42601
rect 23523 42567 23532 42601
rect 23480 42558 23532 42567
rect 23940 42626 23992 42678
rect 24400 42737 24452 42746
rect 24400 42703 24409 42737
rect 24409 42703 24443 42737
rect 24443 42703 24452 42737
rect 24400 42694 24452 42703
rect 24492 42626 24544 42678
rect 26424 42830 26476 42882
rect 28632 42873 28684 42882
rect 28632 42839 28641 42873
rect 28641 42839 28675 42873
rect 28675 42839 28684 42873
rect 28632 42830 28684 42839
rect 29184 42873 29236 42882
rect 29184 42839 29193 42873
rect 29193 42839 29227 42873
rect 29227 42839 29236 42873
rect 29184 42830 29236 42839
rect 29276 42873 29328 42882
rect 29276 42839 29285 42873
rect 29285 42839 29319 42873
rect 29319 42839 29328 42873
rect 29276 42830 29328 42839
rect 30472 42873 30524 42882
rect 30472 42839 30481 42873
rect 30481 42839 30515 42873
rect 30515 42839 30524 42873
rect 30472 42830 30524 42839
rect 30932 42762 30984 42814
rect 27436 42694 27488 42746
rect 26056 42626 26108 42678
rect 26792 42669 26844 42678
rect 26792 42635 26801 42669
rect 26801 42635 26835 42669
rect 26835 42635 26844 42669
rect 26792 42626 26844 42635
rect 28816 42626 28868 42678
rect 29460 42669 29512 42678
rect 29460 42635 29469 42669
rect 29469 42635 29503 42669
rect 29503 42635 29512 42669
rect 29460 42626 29512 42635
rect 30564 42626 30616 42678
rect 25872 42601 25924 42610
rect 25872 42567 25881 42601
rect 25881 42567 25915 42601
rect 25915 42567 25924 42601
rect 25872 42558 25924 42567
rect 8172 42406 8224 42458
rect 8236 42406 8288 42458
rect 8300 42406 8352 42458
rect 8364 42406 8416 42458
rect 8428 42406 8480 42458
rect 15946 42406 15998 42458
rect 16010 42406 16062 42458
rect 16074 42406 16126 42458
rect 16138 42406 16190 42458
rect 16202 42406 16254 42458
rect 23720 42406 23772 42458
rect 23784 42406 23836 42458
rect 23848 42406 23900 42458
rect 23912 42406 23964 42458
rect 23976 42406 24028 42458
rect 31494 42406 31546 42458
rect 31558 42406 31610 42458
rect 31622 42406 31674 42458
rect 31686 42406 31738 42458
rect 31750 42406 31802 42458
rect 11520 42286 11572 42338
rect 12348 42329 12400 42338
rect 12348 42295 12357 42329
rect 12357 42295 12391 42329
rect 12391 42295 12400 42329
rect 12348 42286 12400 42295
rect 12900 42286 12952 42338
rect 13452 42286 13504 42338
rect 13544 42286 13596 42338
rect 13820 42286 13872 42338
rect 14280 42286 14332 42338
rect 14464 42286 14516 42338
rect 2320 42218 2372 42270
rect 3884 42218 3936 42270
rect 11336 42218 11388 42270
rect 12164 42218 12216 42270
rect 3424 42193 3476 42202
rect 3424 42159 3433 42193
rect 3433 42159 3467 42193
rect 3467 42159 3476 42193
rect 3424 42150 3476 42159
rect 12624 42082 12676 42134
rect 13360 42150 13412 42202
rect 14004 42218 14056 42270
rect 14188 42150 14240 42202
rect 14372 42193 14424 42202
rect 14372 42159 14381 42193
rect 14381 42159 14415 42193
rect 14415 42159 14424 42193
rect 14372 42150 14424 42159
rect 15108 42150 15160 42202
rect 15384 42171 15436 42223
rect 15660 42214 15712 42223
rect 15660 42180 15669 42214
rect 15669 42180 15703 42214
rect 15703 42180 15712 42214
rect 15660 42171 15712 42180
rect 16396 42286 16448 42338
rect 16948 42166 17000 42218
rect 17132 42150 17184 42202
rect 17316 42217 17368 42226
rect 17316 42183 17325 42217
rect 17325 42183 17359 42217
rect 17359 42183 17368 42217
rect 17316 42174 17368 42183
rect 17408 42218 17460 42270
rect 19800 42218 19852 42270
rect 22744 42329 22796 42338
rect 22744 42295 22753 42329
rect 22753 42295 22787 42329
rect 22787 42295 22796 42329
rect 22744 42286 22796 42295
rect 23296 42286 23348 42338
rect 24308 42286 24360 42338
rect 1860 42057 1912 42066
rect 1860 42023 1869 42057
rect 1869 42023 1903 42057
rect 1903 42023 1912 42057
rect 1860 42014 1912 42023
rect 4160 42014 4212 42066
rect 11796 42007 11848 42016
rect 11796 41973 11805 42007
rect 11805 41973 11839 42007
rect 11839 41973 11848 42007
rect 11796 41964 11848 41973
rect 11980 42057 12032 42066
rect 11980 42023 11989 42057
rect 11989 42023 12023 42057
rect 12023 42023 12032 42057
rect 11980 42014 12032 42023
rect 12716 42048 12768 42100
rect 15476 42082 15528 42134
rect 15568 42082 15620 42134
rect 12992 42014 13044 42066
rect 13820 42014 13872 42066
rect 14280 42007 14332 42016
rect 14280 41973 14289 42007
rect 14289 41973 14323 42007
rect 14323 41973 14332 42007
rect 14280 41964 14332 41973
rect 14832 42014 14884 42066
rect 16580 42082 16632 42134
rect 16856 42125 16908 42134
rect 16856 42091 16865 42125
rect 16865 42091 16899 42125
rect 16899 42091 16908 42125
rect 16856 42082 16908 42091
rect 19892 42150 19944 42202
rect 20260 42261 20312 42270
rect 20260 42227 20269 42261
rect 20269 42227 20303 42261
rect 20303 42227 20312 42261
rect 20260 42218 20312 42227
rect 20352 42218 20404 42270
rect 21456 42227 21508 42236
rect 21456 42193 21465 42227
rect 21465 42193 21499 42227
rect 21499 42193 21508 42227
rect 21456 42184 21508 42193
rect 21640 42227 21692 42270
rect 21640 42218 21649 42227
rect 21649 42218 21683 42227
rect 21683 42218 21692 42227
rect 21916 42184 21968 42236
rect 22284 42261 22336 42270
rect 22284 42227 22293 42261
rect 22293 42227 22327 42261
rect 22327 42227 22336 42261
rect 22284 42218 22336 42227
rect 22376 42209 22428 42218
rect 22376 42175 22385 42209
rect 22385 42175 22419 42209
rect 22419 42175 22428 42209
rect 22376 42166 22428 42175
rect 22468 42166 22520 42218
rect 24584 42218 24636 42270
rect 18052 42082 18104 42134
rect 19248 42082 19300 42134
rect 19432 42125 19484 42134
rect 19432 42091 19441 42125
rect 19441 42091 19475 42125
rect 19475 42091 19484 42125
rect 19432 42082 19484 42091
rect 23204 42193 23256 42202
rect 23204 42159 23213 42193
rect 23213 42159 23247 42193
rect 23247 42159 23256 42193
rect 23204 42150 23256 42159
rect 24216 42150 24268 42202
rect 25412 42286 25464 42338
rect 25872 42286 25924 42338
rect 20076 42014 20128 42066
rect 20812 42082 20864 42134
rect 21088 42082 21140 42134
rect 21824 42082 21876 42134
rect 20720 42014 20772 42066
rect 20904 42057 20956 42066
rect 20904 42023 20913 42057
rect 20913 42023 20947 42057
rect 20947 42023 20956 42057
rect 20904 42014 20956 42023
rect 21364 42014 21416 42066
rect 22652 42082 22704 42134
rect 22468 42014 22520 42066
rect 25688 42014 25740 42066
rect 206 41862 514 41914
rect 4285 41862 4337 41914
rect 4349 41862 4401 41914
rect 4413 41862 4465 41914
rect 4477 41862 4529 41914
rect 4541 41862 4593 41914
rect 12059 41862 12111 41914
rect 12123 41862 12175 41914
rect 12187 41862 12239 41914
rect 12251 41862 12303 41914
rect 12315 41862 12367 41914
rect 19833 41862 19885 41914
rect 19897 41862 19949 41914
rect 19961 41862 20013 41914
rect 20025 41862 20077 41914
rect 20089 41862 20141 41914
rect 27607 41862 27659 41914
rect 27671 41862 27723 41914
rect 27735 41862 27787 41914
rect 27799 41862 27851 41914
rect 27863 41862 27915 41914
rect 12348 41742 12400 41794
rect 14556 41742 14608 41794
rect 16304 41742 16356 41794
rect 15016 41674 15068 41726
rect 16948 41742 17000 41794
rect 17224 41742 17276 41794
rect 1860 41606 1912 41658
rect 5264 41606 5316 41658
rect 13084 41606 13136 41658
rect 13636 41606 13688 41658
rect 2320 41581 2372 41590
rect 2320 41547 2329 41581
rect 2329 41547 2363 41581
rect 2363 41547 2372 41581
rect 2320 41538 2372 41547
rect 3884 41581 3936 41590
rect 3884 41547 3893 41581
rect 3893 41547 3927 41581
rect 3927 41547 3936 41581
rect 3884 41538 3936 41547
rect 4160 41581 4212 41590
rect 4160 41547 4194 41581
rect 4194 41547 4212 41581
rect 4160 41538 4212 41547
rect 11704 41581 11756 41590
rect 11704 41547 11713 41581
rect 11713 41547 11747 41581
rect 11747 41547 11756 41581
rect 11704 41538 11756 41547
rect 12348 41538 12400 41590
rect 12900 41553 12952 41605
rect 12992 41596 13044 41605
rect 12992 41562 13001 41596
rect 13001 41562 13035 41596
rect 13035 41562 13044 41596
rect 12992 41553 13044 41562
rect 13820 41566 13872 41618
rect 14004 41538 14056 41590
rect 14188 41538 14240 41590
rect 15108 41598 15160 41607
rect 15108 41564 15117 41598
rect 15117 41564 15151 41598
rect 15151 41564 15160 41598
rect 15108 41555 15160 41564
rect 15384 41649 15436 41658
rect 15384 41615 15393 41649
rect 15393 41615 15427 41649
rect 15427 41615 15436 41649
rect 15384 41606 15436 41615
rect 16212 41606 16264 41658
rect 16580 41674 16632 41726
rect 18052 41674 18104 41726
rect 16856 41649 16908 41658
rect 16856 41615 16865 41649
rect 16865 41615 16899 41649
rect 16899 41615 16908 41649
rect 16856 41606 16908 41615
rect 16948 41649 17000 41658
rect 16948 41615 16957 41649
rect 16957 41615 16991 41649
rect 16991 41615 17000 41649
rect 16948 41606 17000 41615
rect 19248 41649 19300 41658
rect 19248 41615 19257 41649
rect 19257 41615 19291 41649
rect 19291 41615 19300 41649
rect 19248 41606 19300 41615
rect 20996 41742 21048 41794
rect 25688 41795 25740 41804
rect 25688 41761 25697 41795
rect 25697 41761 25731 41795
rect 25731 41761 25740 41795
rect 25688 41752 25740 41761
rect 26792 41742 26844 41794
rect 21088 41674 21140 41726
rect 3056 41513 3108 41522
rect 3056 41479 3065 41513
rect 3065 41479 3099 41513
rect 3099 41479 3108 41513
rect 3056 41470 3108 41479
rect 5264 41513 5316 41522
rect 5264 41479 5273 41513
rect 5273 41479 5307 41513
rect 5307 41479 5316 41513
rect 5264 41470 5316 41479
rect 11888 41470 11940 41522
rect 13268 41470 13320 41522
rect 13636 41513 13688 41522
rect 13636 41479 13645 41513
rect 13645 41479 13679 41513
rect 13679 41479 13688 41513
rect 13636 41470 13688 41479
rect 13728 41470 13780 41522
rect 17132 41559 17141 41590
rect 17141 41559 17175 41590
rect 17175 41559 17184 41590
rect 17132 41538 17184 41559
rect 17592 41538 17644 41590
rect 17684 41538 17736 41590
rect 19708 41649 19760 41658
rect 19708 41615 19717 41649
rect 19717 41615 19751 41649
rect 19751 41615 19760 41649
rect 19708 41606 19760 41615
rect 22284 41674 22336 41726
rect 15752 41513 15804 41522
rect 15752 41479 15761 41513
rect 15761 41479 15795 41513
rect 15795 41479 15804 41513
rect 15752 41470 15804 41479
rect 15844 41470 15896 41522
rect 17224 41470 17276 41522
rect 17776 41470 17828 41522
rect 19248 41470 19300 41522
rect 19616 41513 19668 41522
rect 19616 41479 19625 41513
rect 19625 41479 19659 41513
rect 19659 41479 19668 41513
rect 19616 41470 19668 41479
rect 20168 41470 20220 41522
rect 21364 41538 21416 41590
rect 21456 41538 21508 41590
rect 22468 41596 22520 41605
rect 22468 41562 22477 41596
rect 22477 41562 22511 41596
rect 22511 41562 22520 41596
rect 22468 41553 22520 41562
rect 23480 41538 23532 41590
rect 25412 41609 25464 41618
rect 25412 41575 25421 41609
rect 25421 41575 25455 41609
rect 25455 41575 25464 41609
rect 25412 41566 25464 41575
rect 21824 41513 21876 41522
rect 21824 41479 21833 41513
rect 21833 41479 21867 41513
rect 21867 41479 21876 41513
rect 21824 41470 21876 41479
rect 8172 41318 8224 41370
rect 8236 41318 8288 41370
rect 8300 41318 8352 41370
rect 8364 41318 8416 41370
rect 8428 41318 8480 41370
rect 15946 41318 15998 41370
rect 16010 41318 16062 41370
rect 16074 41318 16126 41370
rect 16138 41318 16190 41370
rect 16202 41318 16254 41370
rect 23720 41318 23772 41370
rect 23784 41318 23836 41370
rect 23848 41318 23900 41370
rect 23912 41318 23964 41370
rect 23976 41318 24028 41370
rect 31494 41318 31546 41370
rect 31558 41318 31610 41370
rect 31622 41318 31674 41370
rect 31686 41318 31738 41370
rect 31750 41318 31802 41370
rect 2320 41105 2372 41114
rect 2320 41071 2329 41105
rect 2329 41071 2363 41105
rect 2363 41071 2372 41105
rect 3424 41198 3476 41250
rect 6552 41241 6604 41250
rect 6552 41207 6561 41241
rect 6561 41207 6595 41241
rect 6595 41207 6604 41241
rect 6552 41198 6604 41207
rect 8024 41241 8076 41250
rect 8024 41207 8033 41241
rect 8033 41207 8067 41241
rect 8067 41207 8076 41241
rect 8024 41198 8076 41207
rect 11796 41241 11848 41250
rect 11796 41207 11805 41241
rect 11805 41207 11839 41241
rect 11839 41207 11848 41241
rect 11796 41198 11848 41207
rect 3056 41130 3108 41182
rect 2320 41062 2372 41071
rect 3884 41105 3936 41114
rect 3884 41071 3893 41105
rect 3893 41071 3927 41105
rect 3927 41071 3936 41105
rect 3884 41062 3936 41071
rect 4528 41105 4580 41114
rect 4528 41071 4537 41105
rect 4537 41071 4571 41105
rect 4571 41071 4580 41105
rect 4528 41062 4580 41071
rect 5264 41062 5316 41114
rect 6736 41105 6788 41114
rect 6736 41071 6745 41105
rect 6745 41071 6779 41105
rect 6779 41071 6788 41105
rect 6736 41062 6788 41071
rect 14832 41198 14884 41250
rect 12348 41130 12400 41182
rect 12532 41105 12584 41114
rect 12532 41071 12541 41105
rect 12541 41071 12575 41105
rect 12575 41071 12584 41105
rect 12532 41062 12584 41071
rect 12624 41105 12676 41114
rect 12624 41071 12650 41105
rect 12650 41071 12676 41105
rect 12624 41062 12676 41071
rect 13636 41125 13688 41134
rect 13636 41091 13645 41125
rect 13645 41091 13679 41125
rect 13679 41091 13688 41125
rect 13636 41082 13688 41091
rect 13820 41130 13872 41182
rect 14280 41173 14332 41182
rect 14280 41139 14289 41173
rect 14289 41139 14323 41173
rect 14323 41139 14332 41173
rect 14280 41130 14332 41139
rect 14372 41105 14424 41114
rect 14372 41071 14381 41105
rect 14381 41071 14415 41105
rect 14415 41071 14424 41105
rect 14372 41062 14424 41071
rect 14556 41126 14608 41135
rect 14556 41092 14565 41126
rect 14565 41092 14599 41126
rect 14599 41092 14608 41126
rect 15568 41198 15620 41250
rect 14556 41083 14608 41092
rect 13912 40994 13964 41046
rect 15844 41130 15896 41182
rect 16672 41198 16724 41250
rect 15476 41062 15528 41114
rect 16488 41083 16540 41135
rect 15200 40994 15252 41046
rect 16120 41037 16172 41046
rect 16120 41003 16129 41037
rect 16129 41003 16163 41037
rect 16163 41003 16172 41037
rect 16120 40994 16172 41003
rect 17224 41083 17276 41135
rect 17500 41130 17552 41182
rect 17776 41105 17828 41114
rect 17776 41071 17785 41105
rect 17785 41071 17819 41105
rect 17819 41071 17828 41105
rect 17776 41062 17828 41071
rect 17960 41241 18012 41250
rect 17960 41207 17969 41241
rect 17969 41207 18003 41241
rect 18003 41207 18012 41241
rect 17960 41198 18012 41207
rect 20628 41198 20680 41250
rect 19248 41173 19300 41182
rect 19248 41139 19257 41173
rect 19257 41139 19291 41173
rect 19291 41139 19300 41173
rect 19248 41130 19300 41139
rect 19616 41062 19668 41114
rect 20720 41173 20772 41182
rect 20720 41139 20729 41173
rect 20729 41139 20763 41173
rect 20763 41139 20772 41173
rect 20720 41130 20772 41139
rect 21824 41173 21876 41182
rect 21824 41139 21833 41173
rect 21833 41139 21867 41173
rect 21867 41139 21876 41173
rect 21824 41130 21876 41139
rect 20904 41062 20956 41114
rect 22836 41130 22888 41182
rect 30196 41173 30248 41182
rect 30196 41139 30205 41173
rect 30205 41139 30239 41173
rect 30239 41139 30248 41173
rect 30196 41130 30248 41139
rect 23572 41105 23624 41114
rect 23572 41071 23581 41105
rect 23581 41071 23615 41105
rect 23615 41071 23624 41105
rect 23572 41062 23624 41071
rect 30748 41079 30800 41131
rect 22100 40994 22152 41046
rect 19524 40969 19576 40978
rect 19524 40935 19533 40969
rect 19533 40935 19567 40969
rect 19567 40935 19576 40969
rect 19524 40926 19576 40935
rect 27252 40994 27304 41046
rect 22284 40926 22336 40978
rect 25780 40926 25832 40978
rect 206 40774 514 40826
rect 4285 40774 4337 40826
rect 4349 40774 4401 40826
rect 4413 40774 4465 40826
rect 4477 40774 4529 40826
rect 4541 40774 4593 40826
rect 12059 40774 12111 40826
rect 12123 40774 12175 40826
rect 12187 40774 12239 40826
rect 12251 40774 12303 40826
rect 12315 40774 12367 40826
rect 19833 40774 19885 40826
rect 19897 40774 19949 40826
rect 19961 40774 20013 40826
rect 20025 40774 20077 40826
rect 20089 40774 20141 40826
rect 27607 40774 27659 40826
rect 27671 40774 27723 40826
rect 27735 40774 27787 40826
rect 27799 40774 27851 40826
rect 27863 40774 27915 40826
rect 19524 40654 19576 40706
rect 28724 40654 28776 40706
rect 15384 40586 15436 40638
rect 16948 40586 17000 40638
rect 12440 40450 12492 40502
rect 15200 40508 15252 40517
rect 15200 40474 15209 40508
rect 15209 40474 15243 40508
rect 15243 40474 15252 40508
rect 15200 40465 15252 40474
rect 15660 40508 15712 40517
rect 15660 40474 15669 40508
rect 15669 40474 15703 40508
rect 15703 40474 15712 40508
rect 15660 40465 15712 40474
rect 6736 40382 6788 40434
rect 12808 40382 12860 40434
rect 15752 40450 15804 40502
rect 16948 40382 17000 40434
rect 8172 40230 8224 40282
rect 8236 40230 8288 40282
rect 8300 40230 8352 40282
rect 8364 40230 8416 40282
rect 8428 40230 8480 40282
rect 15946 40230 15998 40282
rect 16010 40230 16062 40282
rect 16074 40230 16126 40282
rect 16138 40230 16190 40282
rect 16202 40230 16254 40282
rect 23720 40230 23772 40282
rect 23784 40230 23836 40282
rect 23848 40230 23900 40282
rect 23912 40230 23964 40282
rect 23976 40230 24028 40282
rect 31494 40230 31546 40282
rect 31558 40230 31610 40282
rect 31622 40230 31674 40282
rect 31686 40230 31738 40282
rect 31750 40230 31802 40282
rect 8148 40040 8502 40048
rect 8148 39976 8502 40040
rect 8148 39968 8502 39976
rect 1058 39740 1150 39792
rect 18212 39738 18300 39790
rect 31530 39494 31760 39752
<< metal2 >>
rect 4526 44822 4582 44831
rect 15842 44822 15898 44831
rect 4526 44757 4582 44766
rect 15752 44786 15804 44792
rect 846 44550 902 44559
rect 846 44485 848 44494
rect 900 44485 902 44494
rect 1582 44550 1638 44559
rect 1582 44485 1584 44494
rect 848 44456 900 44462
rect 1636 44485 1638 44494
rect 2318 44550 2374 44559
rect 2318 44485 2320 44494
rect 1584 44456 1636 44462
rect 2372 44485 2374 44494
rect 3238 44550 3294 44559
rect 3238 44485 3240 44494
rect 2320 44456 2372 44462
rect 3292 44485 3294 44494
rect 3790 44550 3846 44559
rect 4540 44520 4568 44757
rect 15842 44757 15898 44766
rect 17038 44822 17094 44831
rect 25226 44822 25282 44831
rect 17038 44757 17094 44766
rect 23296 44786 23348 44792
rect 15752 44728 15804 44734
rect 9678 44686 9734 44695
rect 8172 44636 8480 44645
rect 8172 44634 8178 44636
rect 8234 44634 8258 44636
rect 8314 44634 8338 44636
rect 8394 44634 8418 44636
rect 8474 44634 8480 44636
rect 8234 44582 8236 44634
rect 8416 44582 8418 44634
rect 9678 44621 9734 44630
rect 8172 44580 8178 44582
rect 8234 44580 8258 44582
rect 8314 44580 8338 44582
rect 8394 44580 8418 44582
rect 8474 44580 8480 44582
rect 8172 44571 8480 44580
rect 5262 44550 5318 44559
rect 3790 44485 3792 44494
rect 3240 44456 3292 44462
rect 3844 44485 3846 44494
rect 4528 44514 4580 44520
rect 3792 44456 3844 44462
rect 5262 44485 5264 44494
rect 4528 44456 4580 44462
rect 5316 44485 5318 44494
rect 5998 44550 6054 44559
rect 5998 44485 6000 44494
rect 5264 44456 5316 44462
rect 6052 44485 6054 44494
rect 6000 44456 6052 44462
rect 9692 44452 9720 44621
rect 14094 44550 14150 44559
rect 13912 44514 13964 44520
rect 14094 44485 14096 44494
rect 13912 44456 13964 44462
rect 14148 44485 14150 44494
rect 15660 44514 15712 44520
rect 14096 44456 14148 44462
rect 15660 44456 15712 44462
rect 9680 44446 9732 44452
rect 13360 44446 13412 44452
rect 9680 44388 9732 44394
rect 12624 44399 12676 44405
rect 13360 44388 13412 44394
rect 13820 44394 13872 44400
rect 12624 44341 12676 44347
rect 12532 44242 12584 44248
rect 12532 44184 12584 44190
rect 206 44092 514 44101
rect 206 44090 212 44092
rect 508 44090 514 44092
rect 206 44036 212 44038
rect 508 44036 514 44038
rect 206 44027 514 44036
rect 4285 44092 4593 44101
rect 4285 44090 4291 44092
rect 4347 44090 4371 44092
rect 4427 44090 4451 44092
rect 4507 44090 4531 44092
rect 4587 44090 4593 44092
rect 4347 44038 4349 44090
rect 4529 44038 4531 44090
rect 4285 44036 4291 44038
rect 4347 44036 4371 44038
rect 4427 44036 4451 44038
rect 4507 44036 4531 44038
rect 4587 44036 4593 44038
rect 4285 44027 4593 44036
rect 12059 44092 12367 44101
rect 12059 44090 12065 44092
rect 12121 44090 12145 44092
rect 12201 44090 12225 44092
rect 12281 44090 12305 44092
rect 12361 44090 12367 44092
rect 12121 44038 12123 44090
rect 12303 44038 12305 44090
rect 12059 44036 12065 44038
rect 12121 44036 12145 44038
rect 12201 44036 12225 44038
rect 12281 44036 12305 44038
rect 12361 44036 12367 44038
rect 12059 44027 12367 44036
rect 11336 43766 11388 43772
rect 11336 43708 11388 43714
rect 11520 43766 11572 43772
rect 11520 43708 11572 43714
rect 11244 43698 11296 43704
rect 11244 43640 11296 43646
rect 8172 43548 8480 43557
rect 8172 43546 8178 43548
rect 8234 43546 8258 43548
rect 8314 43546 8338 43548
rect 8394 43546 8418 43548
rect 8474 43546 8480 43548
rect 8234 43494 8236 43546
rect 8416 43494 8418 43546
rect 8172 43492 8178 43494
rect 8234 43492 8258 43494
rect 8314 43492 8338 43494
rect 8394 43492 8418 43494
rect 8474 43492 8480 43494
rect 8172 43483 8480 43492
rect 206 43004 514 43013
rect 206 43002 212 43004
rect 508 43002 514 43004
rect 206 42948 212 42950
rect 508 42948 514 42950
rect 206 42939 514 42948
rect 4285 43004 4593 43013
rect 4285 43002 4291 43004
rect 4347 43002 4371 43004
rect 4427 43002 4451 43004
rect 4507 43002 4531 43004
rect 4587 43002 4593 43004
rect 4347 42950 4349 43002
rect 4529 42950 4531 43002
rect 4285 42948 4291 42950
rect 4347 42948 4371 42950
rect 4427 42948 4451 42950
rect 4507 42948 4531 42950
rect 4587 42948 4593 42950
rect 4285 42939 4593 42948
rect 11152 42882 11204 42888
rect 11152 42824 11204 42830
rect 11164 42791 11192 42824
rect 11150 42782 11206 42791
rect 11150 42717 11206 42726
rect 8172 42460 8480 42469
rect 8172 42458 8178 42460
rect 8234 42458 8258 42460
rect 8314 42458 8338 42460
rect 8394 42458 8418 42460
rect 8474 42458 8480 42460
rect 8234 42406 8236 42458
rect 8416 42406 8418 42458
rect 8172 42404 8178 42406
rect 8234 42404 8258 42406
rect 8314 42404 8338 42406
rect 8394 42404 8418 42406
rect 8474 42404 8480 42406
rect 8172 42395 8480 42404
rect 2320 42270 2372 42276
rect 2320 42212 2372 42218
rect 3884 42270 3936 42276
rect 11164 42247 11192 42717
rect 3884 42212 3936 42218
rect 11150 42238 11206 42247
rect 1860 42066 1912 42072
rect 1860 42008 1912 42014
rect 206 41916 514 41925
rect 206 41914 212 41916
rect 508 41914 514 41916
rect 206 41860 212 41862
rect 508 41860 514 41862
rect 206 41851 514 41860
rect 1872 41664 1900 42008
rect 1860 41658 1912 41664
rect 1860 41600 1912 41606
rect 2332 41596 2360 42212
rect 3424 42202 3476 42208
rect 3424 42144 3476 42150
rect 2320 41590 2372 41596
rect 2320 41532 2372 41538
rect 3056 41522 3108 41528
rect 3056 41464 3108 41470
rect 3068 41188 3096 41464
rect 3436 41256 3464 42144
rect 3896 41596 3924 42212
rect 11150 42173 11206 42182
rect 11256 42111 11284 43640
rect 11348 43228 11376 43708
rect 11336 43222 11388 43228
rect 11336 43164 11388 43170
rect 11348 42276 11376 43164
rect 11532 42344 11560 43708
rect 11796 43154 11848 43160
rect 11796 43096 11848 43102
rect 11520 42338 11572 42344
rect 11520 42280 11572 42286
rect 11336 42270 11388 42276
rect 11336 42212 11388 42218
rect 11242 42102 11298 42111
rect 4160 42066 4212 42072
rect 11242 42037 11298 42046
rect 11808 42022 11836 43096
rect 12059 43004 12367 43013
rect 12059 43002 12065 43004
rect 12121 43002 12145 43004
rect 12201 43002 12225 43004
rect 12281 43002 12305 43004
rect 12361 43002 12367 43004
rect 12121 42950 12123 43002
rect 12303 42950 12305 43002
rect 12059 42948 12065 42950
rect 12121 42948 12145 42950
rect 12201 42948 12225 42950
rect 12281 42948 12305 42950
rect 12361 42948 12367 42950
rect 12059 42939 12367 42948
rect 12440 42882 12492 42888
rect 12440 42824 12492 42830
rect 11978 42646 12034 42655
rect 11978 42581 12034 42590
rect 12164 42610 12216 42616
rect 11992 42072 12020 42581
rect 12164 42552 12216 42558
rect 12348 42610 12400 42616
rect 12348 42552 12400 42558
rect 12176 42276 12204 42552
rect 12360 42344 12388 42552
rect 12452 42383 12480 42824
rect 12544 42684 12572 44184
rect 12636 43228 12664 44341
rect 13372 44316 13400 44388
rect 13544 44378 13596 44384
rect 13596 44342 13820 44366
rect 13596 44338 13872 44342
rect 13820 44336 13872 44338
rect 13544 44320 13596 44326
rect 13268 44310 13320 44316
rect 13268 44252 13320 44258
rect 13360 44310 13412 44316
rect 13360 44252 13412 44258
rect 13176 44242 13228 44248
rect 13176 44184 13228 44190
rect 13188 43704 13216 44184
rect 13176 43698 13228 43704
rect 13176 43640 13228 43646
rect 13188 43364 13216 43640
rect 13176 43358 13228 43364
rect 13176 43300 13228 43306
rect 13280 43296 13308 44252
rect 13084 43290 13136 43296
rect 13084 43232 13136 43238
rect 13268 43290 13320 43296
rect 13268 43232 13320 43238
rect 12624 43222 12676 43228
rect 12624 43164 12676 43170
rect 12636 42820 12664 43164
rect 13096 42888 13124 43232
rect 13556 43228 13584 44320
rect 13820 44242 13872 44248
rect 13820 44184 13872 44190
rect 13544 43222 13596 43228
rect 13544 43164 13596 43170
rect 13084 42882 13136 42888
rect 13084 42824 13136 42830
rect 12624 42814 12676 42820
rect 12624 42756 12676 42762
rect 13360 42814 13412 42820
rect 13360 42756 13412 42762
rect 12532 42678 12584 42684
rect 12532 42620 12584 42626
rect 12438 42374 12494 42383
rect 12348 42338 12400 42344
rect 12438 42309 12494 42318
rect 12348 42280 12400 42286
rect 12164 42270 12216 42276
rect 12164 42212 12216 42218
rect 11980 42066 12032 42072
rect 4160 42008 4212 42014
rect 11796 42016 11848 42022
rect 4172 41596 4200 42008
rect 11980 42008 12032 42014
rect 11796 41958 11848 41964
rect 4285 41916 4593 41925
rect 4285 41914 4291 41916
rect 4347 41914 4371 41916
rect 4427 41914 4451 41916
rect 4507 41914 4531 41916
rect 4587 41914 4593 41916
rect 4347 41862 4349 41914
rect 4529 41862 4531 41914
rect 4285 41860 4291 41862
rect 4347 41860 4371 41862
rect 4427 41860 4451 41862
rect 4507 41860 4531 41862
rect 4587 41860 4593 41862
rect 4285 41851 4593 41860
rect 12059 41916 12367 41925
rect 12059 41914 12065 41916
rect 12121 41914 12145 41916
rect 12201 41914 12225 41916
rect 12281 41914 12305 41916
rect 12361 41914 12367 41916
rect 12121 41862 12123 41914
rect 12303 41862 12305 41914
rect 12059 41860 12065 41862
rect 12121 41860 12145 41862
rect 12201 41860 12225 41862
rect 12281 41860 12305 41862
rect 12361 41860 12367 41862
rect 12059 41851 12367 41860
rect 11886 41830 11942 41839
rect 11886 41765 11942 41774
rect 12348 41794 12400 41800
rect 5264 41658 5316 41664
rect 5264 41600 5316 41606
rect 3884 41590 3936 41596
rect 3884 41532 3936 41538
rect 4160 41590 4212 41596
rect 4160 41532 4212 41538
rect 3424 41250 3476 41256
rect 3424 41192 3476 41198
rect 3056 41182 3108 41188
rect 2134 41150 2190 41159
rect 3056 41124 3108 41130
rect 3896 41120 3924 41532
rect 5276 41528 5304 41600
rect 11704 41590 11756 41596
rect 11704 41532 11756 41538
rect 5264 41522 5316 41528
rect 5264 41464 5316 41470
rect 4342 41150 4398 41159
rect 2320 41114 2372 41120
rect 2190 41094 2320 41114
rect 2134 41062 2320 41094
rect 2320 41056 2372 41062
rect 3884 41114 3936 41120
rect 5276 41120 5304 41464
rect 8172 41372 8480 41381
rect 8172 41370 8178 41372
rect 8234 41370 8258 41372
rect 8314 41370 8338 41372
rect 8394 41370 8418 41372
rect 8474 41370 8480 41372
rect 8234 41318 8236 41370
rect 8416 41318 8418 41370
rect 8172 41316 8178 41318
rect 8234 41316 8258 41318
rect 8314 41316 8338 41318
rect 8394 41316 8418 41318
rect 8474 41316 8480 41318
rect 8172 41307 8480 41316
rect 11716 41295 11744 41532
rect 11900 41528 11928 41765
rect 12348 41736 12400 41742
rect 12360 41596 12388 41736
rect 12348 41590 12400 41596
rect 12348 41532 12400 41538
rect 11888 41522 11940 41528
rect 11888 41464 11940 41470
rect 11702 41286 11758 41295
rect 6552 41250 6604 41256
rect 6552 41192 6604 41198
rect 8024 41250 8076 41256
rect 11702 41221 11758 41230
rect 11796 41250 11848 41256
rect 8024 41192 8076 41198
rect 11796 41192 11848 41198
rect 6564 41159 6592 41192
rect 8036 41159 8064 41192
rect 11808 41159 11836 41192
rect 12360 41188 12388 41532
rect 12348 41182 12400 41188
rect 6550 41150 6606 41159
rect 4528 41114 4580 41120
rect 4398 41094 4528 41114
rect 4342 41062 4528 41094
rect 3884 41056 3936 41062
rect 4528 41056 4580 41062
rect 5264 41114 5316 41120
rect 8022 41150 8078 41159
rect 6550 41085 6606 41094
rect 6736 41114 6788 41120
rect 5264 41056 5316 41062
rect 8022 41085 8078 41094
rect 11794 41150 11850 41159
rect 12348 41124 12400 41130
rect 11794 41085 11850 41094
rect 6736 41056 6788 41062
rect 206 40828 514 40837
rect 206 40826 212 40828
rect 508 40826 514 40828
rect 206 40772 212 40774
rect 508 40772 514 40774
rect 206 40763 514 40772
rect 4285 40828 4593 40837
rect 4285 40826 4291 40828
rect 4347 40826 4371 40828
rect 4427 40826 4451 40828
rect 4507 40826 4531 40828
rect 4587 40826 4593 40828
rect 4347 40774 4349 40826
rect 4529 40774 4531 40826
rect 4285 40772 4291 40774
rect 4347 40772 4371 40774
rect 4427 40772 4451 40774
rect 4507 40772 4531 40774
rect 4587 40772 4593 40774
rect 4285 40763 4593 40772
rect 6748 40440 6776 41056
rect 12059 40828 12367 40837
rect 12059 40826 12065 40828
rect 12121 40826 12145 40828
rect 12201 40826 12225 40828
rect 12281 40826 12305 40828
rect 12361 40826 12367 40828
rect 12121 40774 12123 40826
rect 12303 40774 12305 40826
rect 12059 40772 12065 40774
rect 12121 40772 12145 40774
rect 12201 40772 12225 40774
rect 12281 40772 12305 40774
rect 12361 40772 12367 40774
rect 12059 40763 12367 40772
rect 12452 40508 12480 42309
rect 12636 42198 12664 42756
rect 12992 42678 13044 42684
rect 12990 42646 12992 42655
rect 13084 42678 13136 42684
rect 13044 42646 13046 42655
rect 13084 42620 13136 42626
rect 12990 42581 13046 42590
rect 12900 42338 12952 42344
rect 12900 42280 12952 42286
rect 12636 42170 12756 42198
rect 12624 42134 12676 42140
rect 12728 42106 12756 42170
rect 12624 42076 12676 42082
rect 12716 42100 12768 42106
rect 12530 41558 12586 41567
rect 12530 41493 12586 41502
rect 12544 41120 12572 41493
rect 12636 41159 12664 42076
rect 12716 42042 12768 42048
rect 12912 41611 12940 42280
rect 12992 42066 13044 42072
rect 12992 42008 13044 42014
rect 13004 41611 13032 42008
rect 13096 41703 13124 42620
rect 13372 42208 13400 42756
rect 13452 42693 13504 42699
rect 13452 42635 13504 42641
rect 13464 42344 13492 42635
rect 13556 42616 13584 43164
rect 13544 42610 13596 42616
rect 13544 42552 13596 42558
rect 13556 42344 13584 42552
rect 13832 42344 13860 44184
rect 13452 42338 13504 42344
rect 13452 42280 13504 42286
rect 13544 42338 13596 42344
rect 13544 42280 13596 42286
rect 13820 42338 13872 42344
rect 13820 42280 13872 42286
rect 13360 42202 13412 42208
rect 13360 42144 13412 42150
rect 13820 42066 13872 42072
rect 13820 42008 13872 42014
rect 13082 41694 13138 41703
rect 13082 41629 13084 41638
rect 12900 41605 12952 41611
rect 12992 41605 13044 41611
rect 12900 41547 12952 41553
rect 12990 41558 12992 41567
rect 13136 41629 13138 41638
rect 13266 41694 13322 41703
rect 13266 41629 13322 41638
rect 13636 41658 13688 41664
rect 13084 41600 13136 41606
rect 13044 41558 13046 41567
rect 13280 41528 13308 41629
rect 13688 41618 13768 41646
rect 13832 41624 13860 42008
rect 13636 41600 13688 41606
rect 13740 41528 13768 41618
rect 13820 41618 13872 41624
rect 13820 41560 13872 41566
rect 12990 41493 13046 41502
rect 13268 41522 13320 41528
rect 13268 41464 13320 41470
rect 13636 41522 13688 41528
rect 13636 41464 13688 41470
rect 13728 41522 13780 41528
rect 13728 41464 13780 41470
rect 12622 41150 12678 41159
rect 12532 41114 12584 41120
rect 13648 41140 13676 41464
rect 13832 41188 13860 41560
rect 13820 41182 13872 41188
rect 12622 41085 12624 41094
rect 12532 41056 12584 41062
rect 12676 41085 12678 41094
rect 13636 41134 13688 41140
rect 13820 41124 13872 41130
rect 13636 41076 13688 41082
rect 12624 41056 12676 41062
rect 13924 41052 13952 44456
rect 14372 44446 14424 44452
rect 14372 44388 14424 44394
rect 14738 44414 14794 44423
rect 14280 44378 14332 44384
rect 14280 44320 14332 44326
rect 14002 43870 14058 43879
rect 14002 43805 14004 43814
rect 14056 43805 14058 43814
rect 14004 43776 14056 43782
rect 14016 43704 14044 43776
rect 14188 43766 14240 43772
rect 14188 43708 14240 43714
rect 14004 43698 14056 43704
rect 14004 43640 14056 43646
rect 14200 43432 14228 43708
rect 14188 43426 14240 43432
rect 14188 43368 14240 43374
rect 14186 43326 14242 43335
rect 14186 43261 14242 43270
rect 14200 42616 14228 43261
rect 14188 42610 14240 42616
rect 14188 42552 14240 42558
rect 14292 42478 14320 44320
rect 14384 43787 14412 44388
rect 14738 44349 14794 44358
rect 15568 44402 15620 44408
rect 14372 43781 14424 43787
rect 14372 43723 14424 43729
rect 14752 43704 14780 44349
rect 15568 44344 15620 44350
rect 14924 44310 14976 44316
rect 14924 44252 14976 44258
rect 15476 44310 15528 44316
rect 15476 44252 15528 44258
rect 14464 43698 14516 43704
rect 14464 43640 14516 43646
rect 14740 43698 14792 43704
rect 14740 43640 14792 43646
rect 14372 43290 14424 43296
rect 14372 43232 14424 43238
rect 14384 42655 14412 43232
rect 14370 42646 14426 42655
rect 14370 42581 14426 42590
rect 14200 42450 14320 42478
rect 14004 42270 14056 42276
rect 14004 42212 14056 42218
rect 14016 41596 14044 42212
rect 14200 42208 14228 42450
rect 14280 42338 14332 42344
rect 14280 42280 14332 42286
rect 14188 42202 14240 42208
rect 14188 42144 14240 42150
rect 14200 41596 14228 42144
rect 14292 42022 14320 42280
rect 14384 42208 14412 42581
rect 14476 42344 14504 43640
rect 14936 43335 14964 44252
rect 15488 43772 15516 44252
rect 15580 43772 15608 44344
rect 15672 44298 15700 44456
rect 15764 44418 15792 44728
rect 15752 44412 15804 44418
rect 15752 44354 15804 44360
rect 15672 44270 15792 44298
rect 15120 43741 15332 43769
rect 14922 43326 14978 43335
rect 14922 43261 14924 43270
rect 14976 43261 14978 43270
rect 14924 43232 14976 43238
rect 14936 42752 14964 43232
rect 14924 42746 14976 42752
rect 14924 42688 14976 42694
rect 15016 42746 15068 42752
rect 15016 42688 15068 42694
rect 14464 42338 14516 42344
rect 14464 42280 14516 42286
rect 14372 42202 14424 42208
rect 14372 42144 14424 42150
rect 14832 42066 14884 42072
rect 14280 42016 14332 42022
rect 14832 42008 14884 42014
rect 14280 41958 14332 41964
rect 14004 41590 14056 41596
rect 14002 41558 14004 41567
rect 14188 41590 14240 41596
rect 14056 41558 14058 41567
rect 14188 41532 14240 41538
rect 14002 41493 14058 41502
rect 14292 41188 14320 41958
rect 14556 41794 14608 41800
rect 14556 41736 14608 41742
rect 14280 41182 14332 41188
rect 14278 41150 14280 41159
rect 14332 41150 14334 41159
rect 14568 41141 14596 41736
rect 14844 41256 14872 42008
rect 15028 41732 15056 42688
rect 15120 42208 15148 43741
rect 15304 43704 15332 43741
rect 15384 43766 15436 43772
rect 15384 43708 15436 43714
rect 15476 43766 15528 43772
rect 15476 43708 15528 43714
rect 15568 43766 15620 43772
rect 15568 43708 15620 43714
rect 15200 43698 15252 43704
rect 15200 43640 15252 43646
rect 15292 43698 15344 43704
rect 15292 43640 15344 43646
rect 15212 43160 15240 43640
rect 15396 43296 15424 43708
rect 15384 43290 15436 43296
rect 15384 43232 15436 43238
rect 15292 43222 15344 43228
rect 15292 43164 15344 43170
rect 15200 43154 15252 43160
rect 15200 43096 15252 43102
rect 15212 42684 15240 43096
rect 15304 42684 15332 43164
rect 15384 42814 15436 42820
rect 15384 42756 15436 42762
rect 15200 42678 15252 42684
rect 15200 42620 15252 42626
rect 15292 42678 15344 42684
rect 15292 42620 15344 42626
rect 15396 42616 15424 42756
rect 15660 42678 15712 42684
rect 15764 42655 15792 44270
rect 15660 42620 15712 42626
rect 15750 42646 15806 42655
rect 15384 42610 15436 42616
rect 15384 42552 15436 42558
rect 15396 42229 15424 42552
rect 15672 42496 15700 42620
rect 15750 42581 15806 42590
rect 15856 42496 15884 44757
rect 15946 44636 16254 44645
rect 15946 44634 15952 44636
rect 16008 44634 16032 44636
rect 16088 44634 16112 44636
rect 16168 44634 16192 44636
rect 16248 44634 16254 44636
rect 16008 44582 16010 44634
rect 16190 44582 16192 44634
rect 15946 44580 15952 44582
rect 16008 44580 16032 44582
rect 16088 44580 16112 44582
rect 16168 44580 16192 44582
rect 16248 44580 16254 44582
rect 15946 44571 16254 44580
rect 17052 44452 17080 44757
rect 23296 44728 23348 44734
rect 23480 44786 23532 44792
rect 25226 44757 25282 44766
rect 30380 44786 30432 44792
rect 23480 44728 23532 44734
rect 17868 44514 17920 44520
rect 19156 44514 19208 44520
rect 17868 44456 17920 44462
rect 18984 44474 19156 44502
rect 17040 44446 17092 44452
rect 16304 44399 16356 44405
rect 16304 44341 16356 44347
rect 16856 44399 16908 44405
rect 17040 44388 17092 44394
rect 17406 44414 17462 44423
rect 16856 44341 16908 44347
rect 17224 44378 17276 44384
rect 15946 43548 16254 43557
rect 15946 43546 15952 43548
rect 16008 43546 16032 43548
rect 16088 43546 16112 43548
rect 16168 43546 16192 43548
rect 16248 43546 16254 43548
rect 16008 43494 16010 43546
rect 16190 43494 16192 43546
rect 15946 43492 15952 43494
rect 16008 43492 16032 43494
rect 16088 43492 16112 43494
rect 16168 43492 16192 43494
rect 16248 43492 16254 43494
rect 15946 43483 16254 43492
rect 16316 43176 16344 44341
rect 16396 44242 16448 44248
rect 16396 44184 16448 44190
rect 16580 44242 16632 44248
rect 16580 44184 16632 44190
rect 16408 43364 16436 44184
rect 16592 43772 16620 44184
rect 16580 43766 16632 43772
rect 16580 43708 16632 43714
rect 16396 43358 16448 43364
rect 16396 43300 16448 43306
rect 16132 43160 16344 43176
rect 16120 43154 16344 43160
rect 16172 43148 16344 43154
rect 16120 43096 16172 43102
rect 16316 42699 16344 43148
rect 16304 42693 16356 42699
rect 16304 42635 16356 42641
rect 15672 42468 15884 42496
rect 15946 42460 16254 42469
rect 15946 42458 15952 42460
rect 16008 42458 16032 42460
rect 16088 42458 16112 42460
rect 16168 42458 16192 42460
rect 16248 42458 16254 42460
rect 16008 42406 16010 42458
rect 16190 42406 16192 42458
rect 15946 42404 15952 42406
rect 16008 42404 16032 42406
rect 16088 42404 16112 42406
rect 16168 42404 16192 42406
rect 16248 42404 16254 42406
rect 15946 42395 16254 42404
rect 16396 42338 16448 42344
rect 16396 42280 16448 42286
rect 15384 42223 15436 42229
rect 15108 42202 15160 42208
rect 15160 42162 15240 42190
rect 15384 42165 15436 42171
rect 15660 42223 15712 42229
rect 15660 42165 15712 42171
rect 15108 42144 15160 42150
rect 15106 41966 15162 41975
rect 15106 41901 15162 41910
rect 15016 41726 15068 41732
rect 15016 41668 15068 41674
rect 15120 41613 15148 41901
rect 15212 41839 15240 42162
rect 15476 42134 15528 42140
rect 15568 42134 15620 42140
rect 15476 42076 15528 42082
rect 15566 42102 15568 42111
rect 15620 42102 15622 42111
rect 15198 41830 15254 41839
rect 15198 41765 15254 41774
rect 15384 41658 15436 41664
rect 15108 41607 15160 41613
rect 15384 41600 15436 41606
rect 15108 41549 15160 41555
rect 14832 41250 14884 41256
rect 14832 41192 14884 41198
rect 14556 41135 14608 41141
rect 14278 41085 14334 41094
rect 14372 41114 14424 41120
rect 14556 41077 14608 41083
rect 14372 41056 14424 41062
rect 13912 41046 13964 41052
rect 13912 40988 13964 40994
rect 12440 40502 12492 40508
rect 12440 40444 12492 40450
rect 6736 40434 6788 40440
rect 6736 40376 6788 40382
rect 12808 40434 12860 40440
rect 12808 40376 12860 40382
rect 8172 40284 8480 40293
rect 8172 40282 8178 40284
rect 8234 40282 8258 40284
rect 8314 40282 8338 40284
rect 8394 40282 8418 40284
rect 8474 40282 8480 40284
rect 8234 40230 8236 40282
rect 8416 40230 8418 40282
rect 8172 40228 8178 40230
rect 8234 40228 8258 40230
rect 8314 40228 8338 40230
rect 8394 40228 8418 40230
rect 8474 40228 8480 40230
rect 8172 40219 8480 40228
rect 12820 40071 12848 40376
rect 14384 40207 14412 41056
rect 15200 41046 15252 41052
rect 15200 40988 15252 40994
rect 15212 40523 15240 40988
rect 15396 40644 15424 41600
rect 15488 41120 15516 42076
rect 15566 42037 15622 42046
rect 15568 41250 15620 41256
rect 15568 41192 15620 41198
rect 15580 41159 15608 41192
rect 15566 41150 15622 41159
rect 15476 41114 15528 41120
rect 15566 41085 15622 41094
rect 15476 41056 15528 41062
rect 15384 40638 15436 40644
rect 15384 40580 15436 40586
rect 15672 40523 15700 42165
rect 16210 42102 16266 42111
rect 16210 42037 16266 42046
rect 16224 41664 16252 42037
rect 16304 41794 16356 41800
rect 16408 41782 16436 42280
rect 16868 42140 16896 44341
rect 17406 44349 17462 44358
rect 17224 44320 17276 44326
rect 17236 43976 17264 44320
rect 17224 43970 17276 43976
rect 17144 43930 17224 43958
rect 17144 43335 17172 43930
rect 17224 43912 17276 43918
rect 17420 43840 17448 44349
rect 17408 43834 17460 43840
rect 17880 43787 17908 44456
rect 18984 44384 19012 44474
rect 19156 44456 19208 44462
rect 19616 44514 19668 44520
rect 19616 44456 19668 44462
rect 19064 44386 19116 44392
rect 18972 44378 19024 44384
rect 19064 44328 19116 44334
rect 19248 44386 19300 44392
rect 19248 44328 19300 44334
rect 18972 44320 19024 44326
rect 19076 43908 19104 44328
rect 19064 43902 19116 43908
rect 19064 43844 19116 43850
rect 17960 43834 18012 43840
rect 17408 43776 17460 43782
rect 17592 43781 17644 43787
rect 17592 43723 17644 43729
rect 17868 43781 17920 43787
rect 17960 43776 18012 43782
rect 17868 43723 17920 43729
rect 17130 43326 17186 43335
rect 17130 43261 17186 43270
rect 17040 43154 17092 43160
rect 16960 43114 17040 43142
rect 16960 42752 16988 43114
rect 17040 43096 17092 43102
rect 17038 42782 17094 42791
rect 16948 42746 17000 42752
rect 17038 42717 17094 42726
rect 16948 42688 17000 42694
rect 16960 42224 16988 42688
rect 16948 42218 17000 42224
rect 16948 42160 17000 42166
rect 16580 42134 16632 42140
rect 16580 42076 16632 42082
rect 16856 42134 16908 42140
rect 16856 42076 16908 42082
rect 16356 41754 16436 41782
rect 16486 41830 16542 41839
rect 16486 41765 16542 41774
rect 16304 41736 16356 41742
rect 16212 41658 16264 41664
rect 16212 41600 16264 41606
rect 15752 41522 15804 41528
rect 15752 41464 15804 41470
rect 15844 41522 15896 41528
rect 15844 41464 15896 41470
rect 15200 40517 15252 40523
rect 15200 40459 15252 40465
rect 15660 40517 15712 40523
rect 15764 40508 15792 41464
rect 15856 41188 15884 41464
rect 15946 41372 16254 41381
rect 15946 41370 15952 41372
rect 16008 41370 16032 41372
rect 16088 41370 16112 41372
rect 16168 41370 16192 41372
rect 16248 41370 16254 41372
rect 16008 41318 16010 41370
rect 16190 41318 16192 41370
rect 15946 41316 15952 41318
rect 16008 41316 16032 41318
rect 16088 41316 16112 41318
rect 16168 41316 16192 41318
rect 16248 41316 16254 41318
rect 15946 41307 16254 41316
rect 15844 41182 15896 41188
rect 15844 41124 15896 41130
rect 16118 41150 16174 41159
rect 16500 41141 16528 41765
rect 16592 41732 16620 42076
rect 16868 41816 16896 42076
rect 16684 41788 16896 41816
rect 16960 41800 16988 42160
rect 16948 41794 17000 41800
rect 16580 41726 16632 41732
rect 16580 41668 16632 41674
rect 16684 41256 16712 41788
rect 16948 41736 17000 41742
rect 16856 41658 16908 41664
rect 16856 41600 16908 41606
rect 16948 41658 17000 41664
rect 16948 41600 17000 41606
rect 16868 41431 16896 41600
rect 16854 41422 16910 41431
rect 16854 41357 16910 41366
rect 16672 41250 16724 41256
rect 16672 41192 16724 41198
rect 16118 41085 16174 41094
rect 16488 41135 16540 41141
rect 16132 41052 16160 41085
rect 16488 41077 16540 41083
rect 16120 41046 16172 41052
rect 16120 40988 16172 40994
rect 16960 40644 16988 41600
rect 17052 41578 17080 42717
rect 17144 42208 17172 43261
rect 17316 43222 17368 43228
rect 17316 43164 17368 43170
rect 17328 42616 17356 43164
rect 17316 42610 17368 42616
rect 17316 42552 17368 42558
rect 17222 42238 17278 42247
rect 17132 42202 17184 42208
rect 17328 42232 17356 42552
rect 17408 42270 17460 42276
rect 17222 42173 17278 42182
rect 17316 42226 17368 42232
rect 17408 42212 17460 42218
rect 17132 42144 17184 42150
rect 17144 42111 17172 42144
rect 17130 42102 17186 42111
rect 17130 42037 17186 42046
rect 17236 41800 17264 42173
rect 17316 42168 17368 42174
rect 17224 41794 17276 41800
rect 17224 41736 17276 41742
rect 17132 41590 17184 41596
rect 17052 41550 17132 41578
rect 17132 41532 17184 41538
rect 17224 41522 17276 41528
rect 17224 41464 17276 41470
rect 17236 41141 17264 41464
rect 17328 41431 17356 42168
rect 17420 41975 17448 42212
rect 17406 41966 17462 41975
rect 17406 41901 17462 41910
rect 17604 41596 17632 43723
rect 17972 43228 18000 43776
rect 18788 43698 18840 43704
rect 18788 43640 18840 43646
rect 18800 43364 18828 43640
rect 19260 43432 19288 44328
rect 19340 44242 19392 44248
rect 19340 44184 19392 44190
rect 19352 43432 19380 44184
rect 19628 43772 19656 44456
rect 21824 44446 21876 44452
rect 21824 44388 21876 44394
rect 21732 44310 21784 44316
rect 21732 44252 21784 44258
rect 21640 44242 21692 44248
rect 21640 44184 21692 44190
rect 19833 44092 20141 44101
rect 19833 44090 19839 44092
rect 19895 44090 19919 44092
rect 19975 44090 19999 44092
rect 20055 44090 20079 44092
rect 20135 44090 20141 44092
rect 19895 44038 19897 44090
rect 20077 44038 20079 44090
rect 19833 44036 19839 44038
rect 19895 44036 19919 44038
rect 19975 44036 19999 44038
rect 20055 44036 20079 44038
rect 20135 44036 20141 44038
rect 19833 44027 20141 44036
rect 19892 43902 19944 43908
rect 19892 43844 19944 43850
rect 19708 43834 19760 43840
rect 19708 43776 19760 43782
rect 19616 43766 19668 43772
rect 19616 43708 19668 43714
rect 19248 43426 19300 43432
rect 19248 43368 19300 43374
rect 19340 43426 19392 43432
rect 19340 43368 19392 43374
rect 19616 43392 19668 43398
rect 18788 43358 18840 43364
rect 18788 43300 18840 43306
rect 19260 43296 19288 43368
rect 19616 43334 19668 43340
rect 19248 43290 19300 43296
rect 19248 43232 19300 43238
rect 17960 43222 18012 43228
rect 17960 43164 18012 43170
rect 19628 42752 19656 43334
rect 19616 42746 19668 42752
rect 19616 42688 19668 42694
rect 18234 42646 18290 42655
rect 18234 42581 18236 42590
rect 18288 42581 18290 42590
rect 18236 42552 18288 42558
rect 18052 42134 18104 42140
rect 18052 42076 18104 42082
rect 19248 42134 19300 42140
rect 19432 42134 19484 42140
rect 19248 42076 19300 42082
rect 19430 42102 19432 42111
rect 19484 42102 19486 42111
rect 18064 41732 18092 42076
rect 18052 41726 18104 41732
rect 18052 41668 18104 41674
rect 19260 41664 19288 42076
rect 19430 42037 19486 42046
rect 19720 41664 19748 43776
rect 19904 43772 19932 43844
rect 21652 43840 21680 44184
rect 21744 44015 21772 44252
rect 21730 44006 21786 44015
rect 21730 43941 21786 43950
rect 21640 43834 21692 43840
rect 21640 43776 21692 43782
rect 19892 43766 19944 43772
rect 19892 43708 19944 43714
rect 19904 43199 19932 43708
rect 21456 43290 21508 43296
rect 21456 43232 21508 43238
rect 19890 43190 19946 43199
rect 19890 43125 19946 43134
rect 19833 43004 20141 43013
rect 19833 43002 19839 43004
rect 19895 43002 19919 43004
rect 19975 43002 19999 43004
rect 20055 43002 20079 43004
rect 20135 43002 20141 43004
rect 19895 42950 19897 43002
rect 20077 42950 20079 43002
rect 19833 42948 19839 42950
rect 19895 42948 19919 42950
rect 19975 42948 19999 42950
rect 20055 42948 20079 42950
rect 20135 42948 20141 42950
rect 19833 42939 20141 42948
rect 21468 42888 21496 43232
rect 21456 42882 21508 42888
rect 21456 42824 21508 42830
rect 20916 42752 21128 42768
rect 20904 42746 21140 42752
rect 20956 42740 21088 42746
rect 20904 42688 20956 42694
rect 21088 42688 21140 42694
rect 19892 42610 19944 42616
rect 19892 42552 19944 42558
rect 20812 42610 20864 42616
rect 20812 42552 20864 42558
rect 21180 42610 21232 42616
rect 21456 42610 21508 42616
rect 21232 42570 21456 42598
rect 21180 42552 21232 42558
rect 21456 42552 21508 42558
rect 19800 42270 19852 42276
rect 19798 42238 19800 42247
rect 19852 42238 19854 42247
rect 19904 42208 19932 42552
rect 20260 42270 20312 42276
rect 20258 42238 20260 42247
rect 20352 42270 20404 42276
rect 20312 42238 20314 42247
rect 19798 42173 19854 42182
rect 19892 42202 19944 42208
rect 20352 42212 20404 42218
rect 20258 42173 20314 42182
rect 19892 42144 19944 42150
rect 20076 42066 20128 42072
rect 20128 42026 20208 42054
rect 20076 42008 20128 42014
rect 19833 41916 20141 41925
rect 19833 41914 19839 41916
rect 19895 41914 19919 41916
rect 19975 41914 19999 41916
rect 20055 41914 20079 41916
rect 20135 41914 20141 41916
rect 19895 41862 19897 41914
rect 20077 41862 20079 41914
rect 19833 41860 19839 41862
rect 19895 41860 19919 41862
rect 19975 41860 19999 41862
rect 20055 41860 20079 41862
rect 20135 41860 20141 41862
rect 19833 41851 20141 41860
rect 19248 41658 19300 41664
rect 19248 41600 19300 41606
rect 19708 41658 19760 41664
rect 19708 41600 19760 41606
rect 17592 41590 17644 41596
rect 17498 41558 17554 41567
rect 17592 41532 17644 41538
rect 17684 41590 17736 41596
rect 17684 41532 17736 41538
rect 17498 41493 17554 41502
rect 17314 41422 17370 41431
rect 17314 41357 17370 41366
rect 17512 41188 17540 41493
rect 17500 41182 17552 41188
rect 17224 41135 17276 41141
rect 17696 41159 17724 41532
rect 20180 41528 20208 42026
rect 20364 41703 20392 42212
rect 20824 42140 20852 42552
rect 20994 42238 21050 42247
rect 21468 42242 21496 42552
rect 21652 42276 21680 43776
rect 21836 42888 21864 44388
rect 21916 44378 21968 44384
rect 22100 44378 22152 44384
rect 21968 44338 22100 44366
rect 21916 44320 21968 44326
rect 22100 44320 22152 44326
rect 23020 44378 23072 44384
rect 23020 44320 23072 44326
rect 23204 44378 23256 44384
rect 23204 44320 23256 44326
rect 21928 43908 21956 44320
rect 22008 44242 22060 44248
rect 22008 44184 22060 44190
rect 22100 44242 22152 44248
rect 22100 44184 22152 44190
rect 22020 43976 22048 44184
rect 22008 43970 22060 43976
rect 22008 43912 22060 43918
rect 21916 43902 21968 43908
rect 21916 43844 21968 43850
rect 21824 42882 21876 42888
rect 21824 42824 21876 42830
rect 21824 42746 21876 42752
rect 21824 42688 21876 42694
rect 21640 42270 21692 42276
rect 20994 42173 21050 42182
rect 21456 42236 21508 42242
rect 21640 42212 21692 42218
rect 21456 42178 21508 42184
rect 20812 42134 20864 42140
rect 20810 42102 20812 42111
rect 20864 42102 20866 42111
rect 20720 42066 20772 42072
rect 20810 42037 20866 42046
rect 20904 42066 20956 42072
rect 20720 42008 20772 42014
rect 20904 42008 20956 42014
rect 20350 41694 20406 41703
rect 20350 41629 20406 41638
rect 17776 41522 17828 41528
rect 17776 41464 17828 41470
rect 19248 41522 19300 41528
rect 19248 41464 19300 41470
rect 19616 41522 19668 41528
rect 19616 41464 19668 41470
rect 20168 41522 20220 41528
rect 20168 41464 20220 41470
rect 17500 41124 17552 41130
rect 17682 41150 17738 41159
rect 17788 41120 17816 41464
rect 17960 41250 18012 41256
rect 17960 41192 18012 41198
rect 17972 41159 18000 41192
rect 19260 41188 19288 41464
rect 19248 41182 19300 41188
rect 17958 41150 18014 41159
rect 17682 41085 17738 41094
rect 17776 41114 17828 41120
rect 17224 41077 17276 41083
rect 19248 41124 19300 41130
rect 19628 41120 19656 41464
rect 20628 41250 20680 41256
rect 20628 41192 20680 41198
rect 20640 41159 20668 41192
rect 20732 41188 20760 42008
rect 20720 41182 20772 41188
rect 20626 41150 20682 41159
rect 17958 41085 18014 41094
rect 19616 41114 19668 41120
rect 17776 41056 17828 41062
rect 20720 41124 20772 41130
rect 20916 41120 20944 42008
rect 21008 41800 21036 42173
rect 21836 42140 21864 42688
rect 21916 42236 21968 42242
rect 22112 42224 22140 44184
rect 22928 43834 22980 43840
rect 22928 43776 22980 43782
rect 22652 43766 22704 43772
rect 22652 43708 22704 43714
rect 22664 43432 22692 43708
rect 22940 43704 22968 43776
rect 23032 43704 23060 44320
rect 23216 43908 23244 44320
rect 23204 43902 23256 43908
rect 23204 43844 23256 43850
rect 23216 43704 23244 43844
rect 22928 43698 22980 43704
rect 22928 43640 22980 43646
rect 23020 43698 23072 43704
rect 23020 43640 23072 43646
rect 23204 43698 23256 43704
rect 23204 43640 23256 43646
rect 22940 43432 22968 43640
rect 22652 43426 22704 43432
rect 22652 43368 22704 43374
rect 22928 43426 22980 43432
rect 22928 43368 22980 43374
rect 22466 43190 22522 43199
rect 22466 43125 22522 43134
rect 22560 43154 22612 43160
rect 22376 42678 22428 42684
rect 22376 42620 22428 42626
rect 21968 42196 22140 42224
rect 22284 42270 22336 42276
rect 22388 42224 22416 42620
rect 22480 42224 22508 43125
rect 22560 43096 22612 43102
rect 22572 42752 22600 43096
rect 22560 42746 22612 42752
rect 22560 42688 22612 42694
rect 22664 42247 22692 43368
rect 23032 42616 23060 43640
rect 23216 43364 23244 43640
rect 23204 43358 23256 43364
rect 23204 43300 23256 43306
rect 23216 42684 23244 43300
rect 23204 42678 23256 42684
rect 23204 42620 23256 42626
rect 22744 42610 22796 42616
rect 22744 42552 22796 42558
rect 23020 42610 23072 42616
rect 23020 42552 23072 42558
rect 22756 42344 22784 42552
rect 22744 42338 22796 42344
rect 22744 42280 22796 42286
rect 22650 42238 22706 42247
rect 22284 42212 22336 42218
rect 22376 42218 22428 42224
rect 21916 42178 21968 42184
rect 21088 42134 21140 42140
rect 21088 42076 21140 42082
rect 21824 42134 21876 42140
rect 21824 42076 21876 42082
rect 20996 41794 21048 41800
rect 20996 41736 21048 41742
rect 21100 41732 21128 42076
rect 21364 42066 21416 42072
rect 21364 42008 21416 42014
rect 21088 41726 21140 41732
rect 21088 41668 21140 41674
rect 21376 41596 21404 42008
rect 22296 41732 22324 42212
rect 22376 42160 22428 42166
rect 22468 42218 22520 42224
rect 23216 42208 23244 42620
rect 23308 42344 23336 44728
rect 23388 43766 23440 43772
rect 23388 43708 23440 43714
rect 23400 43432 23428 43708
rect 23388 43426 23440 43432
rect 23388 43368 23440 43374
rect 23492 42752 23520 44728
rect 23720 44636 24028 44645
rect 23720 44634 23726 44636
rect 23782 44634 23806 44636
rect 23862 44634 23886 44636
rect 23942 44634 23966 44636
rect 24022 44634 24028 44636
rect 23782 44582 23784 44634
rect 23964 44582 23966 44634
rect 23720 44580 23726 44582
rect 23782 44580 23806 44582
rect 23862 44580 23886 44582
rect 23942 44580 23966 44582
rect 24022 44580 24028 44582
rect 23720 44571 24028 44580
rect 25240 44384 25268 44757
rect 30380 44728 30432 44734
rect 25502 44686 25558 44695
rect 25502 44621 25558 44630
rect 26790 44686 26846 44695
rect 26790 44621 26846 44630
rect 28630 44686 28686 44695
rect 28630 44621 28686 44630
rect 25516 44384 25544 44621
rect 26516 44446 26568 44452
rect 26516 44388 26568 44394
rect 25228 44378 25280 44384
rect 25228 44320 25280 44326
rect 25504 44378 25556 44384
rect 25504 44320 25556 44326
rect 24124 44310 24176 44316
rect 24124 44252 24176 44258
rect 26240 44310 26292 44316
rect 26240 44252 26292 44258
rect 23662 44006 23718 44015
rect 23662 43941 23664 43950
rect 23716 43941 23718 43950
rect 23664 43912 23716 43918
rect 23572 43698 23624 43704
rect 23572 43640 23624 43646
rect 23584 43296 23612 43640
rect 23720 43548 24028 43557
rect 23720 43546 23726 43548
rect 23782 43546 23806 43548
rect 23862 43546 23886 43548
rect 23942 43546 23966 43548
rect 24022 43546 24028 43548
rect 23782 43494 23784 43546
rect 23964 43494 23966 43546
rect 23720 43492 23726 43494
rect 23782 43492 23806 43494
rect 23862 43492 23886 43494
rect 23942 43492 23966 43494
rect 24022 43492 24028 43494
rect 23720 43483 24028 43492
rect 23940 43358 23992 43364
rect 23940 43300 23992 43306
rect 23572 43290 23624 43296
rect 23572 43232 23624 43238
rect 23480 42746 23532 42752
rect 23480 42688 23532 42694
rect 23952 42684 23980 43300
rect 24136 42820 24164 44252
rect 24584 43766 24636 43772
rect 24584 43708 24636 43714
rect 24400 43698 24452 43704
rect 24400 43640 24452 43646
rect 24124 42814 24176 42820
rect 24124 42756 24176 42762
rect 24412 42752 24440 43640
rect 24596 43346 24624 43708
rect 25504 43698 25556 43704
rect 25504 43640 25556 43646
rect 25516 43364 25544 43640
rect 24676 43358 24728 43364
rect 24596 43318 24676 43346
rect 24676 43300 24728 43306
rect 25504 43358 25556 43364
rect 25228 43298 25280 43304
rect 25504 43300 25556 43306
rect 25228 43240 25280 43246
rect 25044 43222 25096 43228
rect 24688 43182 25044 43210
rect 24400 42746 24452 42752
rect 24228 42706 24400 42734
rect 23940 42678 23992 42684
rect 23940 42620 23992 42626
rect 23480 42610 23532 42616
rect 23480 42552 23532 42558
rect 23296 42338 23348 42344
rect 23296 42280 23348 42286
rect 22650 42173 22706 42182
rect 23204 42202 23256 42208
rect 22468 42160 22520 42166
rect 22664 42140 22692 42173
rect 23204 42144 23256 42150
rect 22652 42134 22704 42140
rect 22652 42076 22704 42082
rect 22468 42066 22520 42072
rect 22468 42008 22520 42014
rect 22284 41726 22336 41732
rect 22284 41668 22336 41674
rect 22480 41611 22508 42008
rect 22468 41605 22520 41611
rect 21364 41590 21416 41596
rect 21456 41590 21508 41596
rect 21364 41532 21416 41538
rect 21454 41558 21456 41567
rect 21508 41558 21510 41567
rect 23492 41596 23520 42552
rect 23720 42460 24028 42469
rect 23720 42458 23726 42460
rect 23782 42458 23806 42460
rect 23862 42458 23886 42460
rect 23942 42458 23966 42460
rect 24022 42458 24028 42460
rect 23782 42406 23784 42458
rect 23964 42406 23966 42458
rect 23720 42404 23726 42406
rect 23782 42404 23806 42406
rect 23862 42404 23886 42406
rect 23942 42404 23966 42406
rect 24022 42404 24028 42406
rect 23720 42395 24028 42404
rect 24228 42208 24256 42706
rect 24400 42688 24452 42694
rect 24492 42678 24544 42684
rect 24492 42620 24544 42626
rect 24504 42478 24532 42620
rect 24688 42478 24716 43182
rect 25240 43199 25268 43240
rect 26252 43228 26280 44252
rect 26528 43296 26556 44388
rect 26804 44384 26832 44621
rect 28644 44384 28672 44621
rect 30392 44536 30420 44728
rect 31494 44636 31802 44645
rect 31494 44634 31500 44636
rect 31556 44634 31580 44636
rect 31636 44634 31660 44636
rect 31716 44634 31740 44636
rect 31796 44634 31802 44636
rect 31556 44582 31558 44634
rect 31738 44582 31740 44634
rect 31494 44580 31500 44582
rect 31556 44580 31580 44582
rect 31636 44580 31660 44582
rect 31716 44580 31740 44582
rect 31796 44580 31802 44582
rect 31494 44571 31802 44580
rect 30392 44508 30604 44536
rect 26792 44378 26844 44384
rect 26792 44320 26844 44326
rect 27988 44378 28040 44384
rect 27988 44320 28040 44326
rect 28632 44378 28684 44384
rect 28632 44320 28684 44326
rect 27528 44310 27580 44316
rect 27528 44252 27580 44258
rect 26608 44242 26660 44248
rect 26608 44184 26660 44190
rect 27068 44242 27120 44248
rect 27068 44184 27120 44190
rect 26620 43432 26648 44184
rect 26884 43766 26936 43772
rect 26884 43708 26936 43714
rect 26896 43432 26924 43708
rect 26608 43426 26660 43432
rect 26608 43368 26660 43374
rect 26884 43426 26936 43432
rect 26884 43368 26936 43374
rect 27080 43296 27108 44184
rect 27540 43976 27568 44252
rect 27607 44092 27915 44101
rect 27607 44090 27613 44092
rect 27669 44090 27693 44092
rect 27749 44090 27773 44092
rect 27829 44090 27853 44092
rect 27909 44090 27915 44092
rect 27669 44038 27671 44090
rect 27851 44038 27853 44090
rect 27607 44036 27613 44038
rect 27669 44036 27693 44038
rect 27749 44036 27773 44038
rect 27829 44036 27853 44038
rect 27909 44036 27915 44038
rect 27607 44027 27915 44036
rect 27528 43970 27580 43976
rect 27528 43912 27580 43918
rect 28000 43704 28028 44320
rect 29184 44310 29236 44316
rect 29184 44252 29236 44258
rect 28078 44142 28134 44151
rect 28078 44077 28134 44086
rect 28092 43976 28120 44077
rect 28080 43970 28132 43976
rect 28080 43912 28132 43918
rect 28908 43970 28960 43976
rect 28908 43912 28960 43918
rect 28814 43870 28870 43879
rect 28814 43805 28870 43814
rect 27988 43698 28040 43704
rect 27988 43640 28040 43646
rect 28356 43698 28408 43704
rect 28356 43640 28408 43646
rect 28632 43698 28684 43704
rect 28632 43640 28684 43646
rect 28000 43364 28028 43640
rect 28368 43432 28396 43640
rect 28356 43426 28408 43432
rect 28356 43368 28408 43374
rect 27988 43358 28040 43364
rect 27988 43300 28040 43306
rect 26516 43290 26568 43296
rect 26516 43232 26568 43238
rect 27068 43290 27120 43296
rect 27068 43232 27120 43238
rect 26056 43222 26108 43228
rect 25044 43164 25096 43170
rect 25226 43190 25282 43199
rect 25226 43125 25282 43134
rect 26054 43190 26056 43199
rect 26240 43222 26292 43228
rect 26108 43190 26110 43199
rect 26240 43164 26292 43170
rect 27436 43222 27488 43228
rect 27436 43164 27488 43170
rect 26054 43125 26110 43134
rect 26424 43154 26476 43160
rect 26068 42684 26096 43125
rect 26424 43096 26476 43102
rect 26436 42888 26464 43096
rect 26424 42882 26476 42888
rect 26424 42824 26476 42830
rect 27448 42752 27476 43164
rect 27607 43004 27915 43013
rect 27607 43002 27613 43004
rect 27669 43002 27693 43004
rect 27749 43002 27773 43004
rect 27829 43002 27853 43004
rect 27909 43002 27915 43004
rect 27669 42950 27671 43002
rect 27851 42950 27853 43002
rect 27607 42948 27613 42950
rect 27669 42948 27693 42950
rect 27749 42948 27773 42950
rect 27829 42948 27853 42950
rect 27909 42948 27915 42950
rect 27607 42939 27915 42948
rect 28644 42888 28672 43640
rect 28632 42882 28684 42888
rect 28632 42824 28684 42830
rect 27436 42746 27488 42752
rect 27436 42688 27488 42694
rect 28828 42684 28856 43805
rect 28920 43296 28948 43912
rect 29000 43766 29052 43772
rect 29000 43708 29052 43714
rect 28908 43290 28960 43296
rect 28908 43232 28960 43238
rect 29012 43228 29040 43708
rect 29000 43222 29052 43228
rect 29000 43164 29052 43170
rect 29196 42888 29224 44252
rect 29460 44242 29512 44248
rect 29460 44184 29512 44190
rect 29276 43766 29328 43772
rect 29276 43708 29328 43714
rect 29288 42888 29316 43708
rect 29368 43698 29420 43704
rect 29368 43640 29420 43646
rect 29380 43296 29408 43640
rect 29368 43290 29420 43296
rect 29368 43232 29420 43238
rect 29184 42882 29236 42888
rect 29184 42824 29236 42830
rect 29276 42882 29328 42888
rect 29276 42824 29328 42830
rect 29472 42684 29500 44184
rect 29550 44142 29606 44151
rect 29550 44077 29606 44086
rect 29564 43432 29592 44077
rect 30392 43976 30420 44508
rect 30576 44384 30604 44508
rect 31116 44514 31168 44520
rect 31116 44456 31168 44462
rect 30472 44378 30524 44384
rect 30472 44320 30524 44326
rect 30564 44378 30616 44384
rect 30564 44320 30616 44326
rect 30484 43976 30512 44320
rect 30840 44310 30892 44316
rect 30840 44252 30892 44258
rect 30564 44242 30616 44248
rect 30564 44184 30616 44190
rect 30380 43970 30432 43976
rect 30380 43912 30432 43918
rect 30472 43970 30524 43976
rect 30472 43912 30524 43918
rect 29552 43426 29604 43432
rect 29552 43368 29604 43374
rect 30472 43358 30524 43364
rect 30472 43300 30524 43306
rect 30484 42888 30512 43300
rect 30472 42882 30524 42888
rect 30472 42824 30524 42830
rect 30576 42684 30604 44184
rect 30852 43432 30880 44252
rect 30930 44006 30986 44015
rect 30930 43941 30986 43950
rect 30840 43426 30892 43432
rect 30840 43368 30892 43374
rect 30944 42820 30972 43941
rect 31128 43840 31156 44456
rect 31116 43834 31168 43840
rect 31116 43776 31168 43782
rect 31128 43160 31156 43776
rect 31494 43548 31802 43557
rect 31494 43546 31500 43548
rect 31556 43546 31580 43548
rect 31636 43546 31660 43548
rect 31716 43546 31740 43548
rect 31796 43546 31802 43548
rect 31556 43494 31558 43546
rect 31738 43494 31740 43546
rect 31494 43492 31500 43494
rect 31556 43492 31580 43494
rect 31636 43492 31660 43494
rect 31716 43492 31740 43494
rect 31796 43492 31802 43494
rect 31494 43483 31802 43492
rect 31116 43154 31168 43160
rect 31116 43096 31168 43102
rect 30932 42814 30984 42820
rect 30932 42756 30984 42762
rect 26056 42678 26108 42684
rect 26056 42620 26108 42626
rect 26792 42678 26844 42684
rect 26792 42620 26844 42626
rect 28816 42678 28868 42684
rect 28816 42620 28868 42626
rect 29460 42678 29512 42684
rect 29460 42620 29512 42626
rect 30564 42678 30616 42684
rect 30564 42620 30616 42626
rect 25872 42610 25924 42616
rect 25872 42552 25924 42558
rect 24320 42450 24532 42478
rect 24596 42450 24716 42478
rect 24320 42344 24348 42450
rect 24308 42338 24360 42344
rect 24308 42280 24360 42286
rect 24596 42276 24624 42450
rect 25884 42344 25912 42552
rect 25412 42338 25464 42344
rect 25412 42280 25464 42286
rect 25872 42338 25924 42344
rect 25872 42280 25924 42286
rect 24584 42270 24636 42276
rect 24584 42212 24636 42218
rect 24216 42202 24268 42208
rect 24216 42144 24268 42150
rect 25424 41624 25452 42280
rect 25688 42066 25740 42072
rect 25688 42008 25740 42014
rect 25700 41810 25728 42008
rect 25688 41804 25740 41810
rect 26804 41800 26832 42620
rect 31494 42460 31802 42469
rect 31494 42458 31500 42460
rect 31556 42458 31580 42460
rect 31636 42458 31660 42460
rect 31716 42458 31740 42460
rect 31796 42458 31802 42460
rect 31556 42406 31558 42458
rect 31738 42406 31740 42458
rect 31494 42404 31500 42406
rect 31556 42404 31580 42406
rect 31636 42404 31660 42406
rect 31716 42404 31740 42406
rect 31796 42404 31802 42406
rect 31494 42395 31802 42404
rect 27607 41916 27915 41925
rect 27607 41914 27613 41916
rect 27669 41914 27693 41916
rect 27749 41914 27773 41916
rect 27829 41914 27853 41916
rect 27909 41914 27915 41916
rect 27669 41862 27671 41914
rect 27851 41862 27853 41914
rect 27607 41860 27613 41862
rect 27669 41860 27693 41862
rect 27749 41860 27773 41862
rect 27829 41860 27853 41862
rect 27909 41860 27915 41862
rect 27607 41851 27915 41860
rect 30746 41830 30802 41839
rect 25688 41746 25740 41752
rect 26792 41794 26844 41800
rect 30746 41765 30802 41774
rect 26792 41736 26844 41742
rect 25412 41618 25464 41624
rect 22468 41547 22520 41553
rect 23480 41590 23532 41596
rect 25412 41560 25464 41566
rect 23480 41532 23532 41538
rect 21454 41493 21510 41502
rect 21824 41522 21876 41528
rect 21824 41464 21876 41470
rect 21836 41188 21864 41464
rect 23720 41372 24028 41381
rect 23720 41370 23726 41372
rect 23782 41370 23806 41372
rect 23862 41370 23886 41372
rect 23942 41370 23966 41372
rect 24022 41370 24028 41372
rect 23782 41318 23784 41370
rect 23964 41318 23966 41370
rect 23720 41316 23726 41318
rect 23782 41316 23806 41318
rect 23862 41316 23886 41318
rect 23942 41316 23966 41318
rect 24022 41316 24028 41318
rect 23720 41307 24028 41316
rect 21824 41182 21876 41188
rect 22836 41182 22888 41188
rect 21824 41124 21876 41130
rect 22834 41150 22836 41159
rect 30196 41182 30248 41188
rect 22888 41150 22890 41159
rect 20626 41085 20682 41094
rect 20904 41114 20956 41120
rect 19616 41056 19668 41062
rect 22834 41085 22890 41094
rect 23570 41150 23626 41159
rect 23570 41085 23572 41094
rect 20904 41056 20956 41062
rect 23624 41085 23626 41094
rect 25778 41150 25834 41159
rect 25778 41085 25834 41094
rect 30194 41150 30196 41159
rect 30248 41150 30250 41159
rect 30760 41137 30788 41765
rect 31494 41372 31802 41381
rect 31494 41370 31500 41372
rect 31556 41370 31580 41372
rect 31636 41370 31660 41372
rect 31716 41370 31740 41372
rect 31796 41370 31802 41372
rect 31556 41318 31558 41370
rect 31738 41318 31740 41370
rect 31494 41316 31500 41318
rect 31556 41316 31580 41318
rect 31636 41316 31660 41318
rect 31716 41316 31740 41318
rect 31796 41316 31802 41318
rect 31494 41307 31802 41316
rect 30194 41085 30250 41094
rect 30748 41131 30800 41137
rect 23572 41056 23624 41062
rect 22100 41046 22152 41052
rect 22152 40994 22324 41000
rect 22100 40988 22324 40994
rect 22112 40984 22324 40988
rect 25792 40984 25820 41085
rect 30748 41073 30800 41079
rect 27252 41046 27304 41052
rect 27252 40988 27304 40994
rect 19524 40978 19576 40984
rect 22112 40978 22336 40984
rect 22112 40972 22284 40978
rect 19524 40920 19576 40926
rect 22284 40920 22336 40926
rect 25780 40978 25832 40984
rect 25780 40920 25832 40926
rect 19536 40712 19564 40920
rect 19833 40828 20141 40837
rect 19833 40826 19839 40828
rect 19895 40826 19919 40828
rect 19975 40826 19999 40828
rect 20055 40826 20079 40828
rect 20135 40826 20141 40828
rect 19895 40774 19897 40826
rect 20077 40774 20079 40826
rect 19833 40772 19839 40774
rect 19895 40772 19919 40774
rect 19975 40772 19999 40774
rect 20055 40772 20079 40774
rect 20135 40772 20141 40774
rect 19833 40763 20141 40772
rect 19524 40706 19576 40712
rect 19524 40648 19576 40654
rect 16948 40638 17000 40644
rect 16948 40580 17000 40586
rect 15660 40459 15712 40465
rect 15752 40502 15804 40508
rect 15752 40444 15804 40450
rect 16948 40434 17000 40440
rect 16948 40376 17000 40382
rect 15946 40284 16254 40293
rect 15946 40282 15952 40284
rect 16008 40282 16032 40284
rect 16088 40282 16112 40284
rect 16168 40282 16192 40284
rect 16248 40282 16254 40284
rect 16008 40230 16010 40282
rect 16190 40230 16192 40282
rect 15946 40228 15952 40230
rect 16008 40228 16032 40230
rect 16088 40228 16112 40230
rect 16168 40228 16192 40230
rect 16248 40228 16254 40230
rect 15946 40219 16254 40228
rect 14370 40198 14426 40207
rect 14370 40133 14426 40142
rect 16960 40071 16988 40376
rect 27264 40343 27292 40988
rect 27607 40828 27915 40837
rect 27607 40826 27613 40828
rect 27669 40826 27693 40828
rect 27749 40826 27773 40828
rect 27829 40826 27853 40828
rect 27909 40826 27915 40828
rect 27669 40774 27671 40826
rect 27851 40774 27853 40826
rect 27607 40772 27613 40774
rect 27669 40772 27693 40774
rect 27749 40772 27773 40774
rect 27829 40772 27853 40774
rect 27909 40772 27915 40774
rect 27607 40763 27915 40772
rect 28724 40706 28776 40712
rect 28724 40648 28776 40654
rect 27250 40334 27306 40343
rect 23720 40284 24028 40293
rect 23720 40282 23726 40284
rect 23782 40282 23806 40284
rect 23862 40282 23886 40284
rect 23942 40282 23966 40284
rect 24022 40282 24028 40284
rect 23782 40230 23784 40282
rect 23964 40230 23966 40282
rect 27250 40269 27306 40278
rect 23720 40228 23726 40230
rect 23782 40228 23806 40230
rect 23862 40228 23886 40230
rect 23942 40228 23966 40230
rect 24022 40228 24028 40230
rect 23720 40219 24028 40228
rect 28736 40207 28764 40648
rect 31494 40284 31802 40293
rect 31494 40282 31500 40284
rect 31556 40282 31580 40284
rect 31636 40282 31660 40284
rect 31716 40282 31740 40284
rect 31796 40282 31802 40284
rect 31556 40230 31558 40282
rect 31738 40230 31740 40282
rect 31494 40228 31500 40230
rect 31556 40228 31580 40230
rect 31636 40228 31660 40230
rect 31716 40228 31740 40230
rect 31796 40228 31802 40230
rect 31494 40219 31802 40228
rect 28722 40198 28778 40207
rect 28722 40133 28778 40142
rect 12806 40062 12862 40071
rect 8128 40048 8522 40054
rect 8128 39968 8148 40048
rect 8502 39968 8522 40048
rect 12806 39997 12862 40006
rect 16946 40062 17002 40071
rect 16946 39997 17002 40006
rect 8128 39962 8522 39968
rect 8860 39896 10470 39968
rect 1050 39792 1158 39802
rect 1050 39736 1058 39792
rect 1150 39736 1158 39792
rect 1050 39726 1158 39736
rect 2972 39800 3080 39802
rect 8860 39800 8930 39896
rect 2972 39792 8930 39800
rect 2972 39736 2980 39792
rect 3072 39736 8930 39792
rect 2972 39728 8930 39736
rect 10400 39800 10470 39896
rect 18202 39800 18310 39802
rect 10400 39790 18310 39800
rect 10400 39738 18212 39790
rect 18300 39738 18310 39790
rect 10400 39728 18310 39738
rect 2972 39726 3080 39728
rect 18202 39726 18310 39728
rect 31514 39752 31776 39764
rect 534 39662 608 39672
rect 534 39606 542 39662
rect 598 39606 608 39662
rect 534 39598 608 39606
rect 31400 39662 31474 39672
rect 31400 39606 31410 39662
rect 31466 39606 31474 39662
rect 31400 39598 31474 39606
rect 534 33296 567 39598
rect 599 39530 673 39540
rect 599 39474 607 39530
rect 663 39474 673 39530
rect 599 39466 673 39474
rect 31335 39530 31409 39540
rect 31335 39474 31345 39530
rect 31401 39474 31409 39530
rect 31335 39466 31409 39474
rect 599 33296 632 39466
rect 664 39398 738 39408
rect 664 39342 672 39398
rect 728 39342 738 39398
rect 664 39334 738 39342
rect 31270 39398 31344 39408
rect 31270 39342 31280 39398
rect 31336 39342 31344 39398
rect 31270 39334 31344 39342
rect 664 33296 697 39334
rect 729 39266 803 39276
rect 729 39210 737 39266
rect 793 39210 803 39266
rect 729 39202 803 39210
rect 31205 39266 31279 39276
rect 31205 39210 31215 39266
rect 31271 39210 31279 39266
rect 31205 39202 31279 39210
rect 729 33296 762 39202
rect 794 39134 868 39144
rect 794 39078 802 39134
rect 858 39078 868 39134
rect 794 39070 868 39078
rect 31140 39134 31214 39144
rect 31140 39078 31150 39134
rect 31206 39078 31214 39134
rect 31140 39070 31214 39078
rect 794 33296 827 39070
rect 859 39002 933 39012
rect 859 38946 867 39002
rect 923 38946 933 39002
rect 859 38938 933 38946
rect 31075 39002 31149 39012
rect 31075 38946 31085 39002
rect 31141 38946 31149 39002
rect 31075 38938 31149 38946
rect 859 33296 892 38938
rect 924 38870 998 38880
rect 924 38814 932 38870
rect 988 38814 998 38870
rect 924 38806 998 38814
rect 31010 38870 31084 38880
rect 31010 38814 31020 38870
rect 31076 38814 31084 38870
rect 31010 38806 31084 38814
rect 924 33296 957 38806
rect 989 38738 1063 38748
rect 989 38682 997 38738
rect 1053 38682 1063 38738
rect 989 38674 1063 38682
rect 30945 38738 31019 38748
rect 30945 38682 30955 38738
rect 31011 38682 31019 38738
rect 30945 38674 31019 38682
rect 989 33296 1022 38674
rect 1054 38606 1128 38616
rect 1054 38550 1062 38606
rect 1118 38550 1128 38606
rect 1054 38542 1128 38550
rect 30880 38606 30954 38616
rect 30880 38550 30890 38606
rect 30946 38550 30954 38606
rect 30880 38542 30954 38550
rect 1054 33296 1087 38542
rect 1119 38474 1193 38484
rect 1119 38418 1127 38474
rect 1183 38418 1193 38474
rect 1119 38410 1193 38418
rect 30815 38474 30889 38484
rect 30815 38418 30825 38474
rect 30881 38418 30889 38474
rect 30815 38410 30889 38418
rect 1119 33296 1152 38410
rect 1184 38342 1258 38352
rect 1184 38286 1192 38342
rect 1248 38286 1258 38342
rect 1184 38278 1258 38286
rect 30750 38342 30824 38352
rect 30750 38286 30760 38342
rect 30816 38286 30824 38342
rect 30750 38278 30824 38286
rect 1184 33296 1217 38278
rect 1249 38210 1323 38220
rect 1249 38154 1257 38210
rect 1313 38154 1323 38210
rect 1249 38146 1323 38154
rect 30685 38210 30759 38220
rect 30685 38154 30695 38210
rect 30751 38154 30759 38210
rect 30685 38146 30759 38154
rect 1249 33296 1282 38146
rect 1314 38078 1388 38088
rect 1314 38022 1322 38078
rect 1378 38022 1388 38078
rect 1314 38014 1388 38022
rect 30620 38078 30694 38088
rect 30620 38022 30630 38078
rect 30686 38022 30694 38078
rect 30620 38014 30694 38022
rect 1314 33296 1347 38014
rect 1379 37946 1453 37956
rect 1379 37890 1387 37946
rect 1443 37890 1453 37946
rect 1379 37882 1453 37890
rect 30555 37946 30629 37956
rect 30555 37890 30565 37946
rect 30621 37890 30629 37946
rect 30555 37882 30629 37890
rect 1379 33296 1412 37882
rect 1444 37814 1518 37824
rect 1444 37758 1452 37814
rect 1508 37758 1518 37814
rect 1444 37750 1518 37758
rect 30490 37814 30564 37824
rect 30490 37758 30500 37814
rect 30556 37758 30564 37814
rect 30490 37750 30564 37758
rect 1444 33296 1477 37750
rect 1509 37682 1583 37692
rect 1509 37626 1517 37682
rect 1573 37626 1583 37682
rect 1509 37618 1583 37626
rect 30425 37682 30499 37692
rect 30425 37626 30435 37682
rect 30491 37626 30499 37682
rect 30425 37618 30499 37626
rect 1509 33296 1542 37618
rect 1574 37550 1648 37560
rect 1574 37494 1582 37550
rect 1638 37494 1648 37550
rect 1574 37486 1648 37494
rect 30360 37550 30434 37560
rect 30360 37494 30370 37550
rect 30426 37494 30434 37550
rect 30360 37486 30434 37494
rect 1574 33296 1607 37486
rect 30401 33296 30434 37486
rect 30466 33296 30499 37618
rect 30531 33296 30564 37750
rect 30596 33296 30629 37882
rect 30661 33296 30694 38014
rect 30726 33296 30759 38146
rect 30791 33296 30824 38278
rect 30856 33296 30889 38410
rect 30921 33296 30954 38542
rect 30986 33296 31019 38674
rect 31051 33296 31084 38806
rect 31116 33296 31149 38938
rect 31181 33296 31214 39070
rect 31246 33296 31279 39202
rect 31311 33296 31344 39334
rect 31376 33176 31409 39466
rect 31441 29510 31474 39598
rect 31514 39494 31530 39752
rect 31764 39494 31776 39752
rect 31514 39482 31776 39494
<< via2 >>
rect 4526 44766 4582 44822
rect 846 44514 902 44550
rect 846 44494 848 44514
rect 848 44494 900 44514
rect 900 44494 902 44514
rect 1582 44514 1638 44550
rect 1582 44494 1584 44514
rect 1584 44494 1636 44514
rect 1636 44494 1638 44514
rect 2318 44514 2374 44550
rect 2318 44494 2320 44514
rect 2320 44494 2372 44514
rect 2372 44494 2374 44514
rect 3238 44514 3294 44550
rect 3238 44494 3240 44514
rect 3240 44494 3292 44514
rect 3292 44494 3294 44514
rect 3790 44514 3846 44550
rect 15842 44766 15898 44822
rect 17038 44766 17094 44822
rect 8178 44634 8234 44636
rect 8258 44634 8314 44636
rect 8338 44634 8394 44636
rect 8418 44634 8474 44636
rect 8178 44582 8224 44634
rect 8224 44582 8234 44634
rect 8258 44582 8288 44634
rect 8288 44582 8300 44634
rect 8300 44582 8314 44634
rect 8338 44582 8352 44634
rect 8352 44582 8364 44634
rect 8364 44582 8394 44634
rect 8418 44582 8428 44634
rect 8428 44582 8474 44634
rect 9678 44630 9734 44686
rect 8178 44580 8234 44582
rect 8258 44580 8314 44582
rect 8338 44580 8394 44582
rect 8418 44580 8474 44582
rect 3790 44494 3792 44514
rect 3792 44494 3844 44514
rect 3844 44494 3846 44514
rect 5262 44514 5318 44550
rect 5262 44494 5264 44514
rect 5264 44494 5316 44514
rect 5316 44494 5318 44514
rect 5998 44514 6054 44550
rect 5998 44494 6000 44514
rect 6000 44494 6052 44514
rect 6052 44494 6054 44514
rect 14094 44514 14150 44550
rect 14094 44494 14096 44514
rect 14096 44494 14148 44514
rect 14148 44494 14150 44514
rect 212 44090 508 44092
rect 212 44038 508 44090
rect 212 44036 508 44038
rect 4291 44090 4347 44092
rect 4371 44090 4427 44092
rect 4451 44090 4507 44092
rect 4531 44090 4587 44092
rect 4291 44038 4337 44090
rect 4337 44038 4347 44090
rect 4371 44038 4401 44090
rect 4401 44038 4413 44090
rect 4413 44038 4427 44090
rect 4451 44038 4465 44090
rect 4465 44038 4477 44090
rect 4477 44038 4507 44090
rect 4531 44038 4541 44090
rect 4541 44038 4587 44090
rect 4291 44036 4347 44038
rect 4371 44036 4427 44038
rect 4451 44036 4507 44038
rect 4531 44036 4587 44038
rect 12065 44090 12121 44092
rect 12145 44090 12201 44092
rect 12225 44090 12281 44092
rect 12305 44090 12361 44092
rect 12065 44038 12111 44090
rect 12111 44038 12121 44090
rect 12145 44038 12175 44090
rect 12175 44038 12187 44090
rect 12187 44038 12201 44090
rect 12225 44038 12239 44090
rect 12239 44038 12251 44090
rect 12251 44038 12281 44090
rect 12305 44038 12315 44090
rect 12315 44038 12361 44090
rect 12065 44036 12121 44038
rect 12145 44036 12201 44038
rect 12225 44036 12281 44038
rect 12305 44036 12361 44038
rect 8178 43546 8234 43548
rect 8258 43546 8314 43548
rect 8338 43546 8394 43548
rect 8418 43546 8474 43548
rect 8178 43494 8224 43546
rect 8224 43494 8234 43546
rect 8258 43494 8288 43546
rect 8288 43494 8300 43546
rect 8300 43494 8314 43546
rect 8338 43494 8352 43546
rect 8352 43494 8364 43546
rect 8364 43494 8394 43546
rect 8418 43494 8428 43546
rect 8428 43494 8474 43546
rect 8178 43492 8234 43494
rect 8258 43492 8314 43494
rect 8338 43492 8394 43494
rect 8418 43492 8474 43494
rect 212 43002 508 43004
rect 212 42950 508 43002
rect 212 42948 508 42950
rect 4291 43002 4347 43004
rect 4371 43002 4427 43004
rect 4451 43002 4507 43004
rect 4531 43002 4587 43004
rect 4291 42950 4337 43002
rect 4337 42950 4347 43002
rect 4371 42950 4401 43002
rect 4401 42950 4413 43002
rect 4413 42950 4427 43002
rect 4451 42950 4465 43002
rect 4465 42950 4477 43002
rect 4477 42950 4507 43002
rect 4531 42950 4541 43002
rect 4541 42950 4587 43002
rect 4291 42948 4347 42950
rect 4371 42948 4427 42950
rect 4451 42948 4507 42950
rect 4531 42948 4587 42950
rect 11150 42726 11206 42782
rect 8178 42458 8234 42460
rect 8258 42458 8314 42460
rect 8338 42458 8394 42460
rect 8418 42458 8474 42460
rect 8178 42406 8224 42458
rect 8224 42406 8234 42458
rect 8258 42406 8288 42458
rect 8288 42406 8300 42458
rect 8300 42406 8314 42458
rect 8338 42406 8352 42458
rect 8352 42406 8364 42458
rect 8364 42406 8394 42458
rect 8418 42406 8428 42458
rect 8428 42406 8474 42458
rect 8178 42404 8234 42406
rect 8258 42404 8314 42406
rect 8338 42404 8394 42406
rect 8418 42404 8474 42406
rect 212 41914 508 41916
rect 212 41862 508 41914
rect 212 41860 508 41862
rect 11150 42182 11206 42238
rect 11242 42046 11298 42102
rect 12065 43002 12121 43004
rect 12145 43002 12201 43004
rect 12225 43002 12281 43004
rect 12305 43002 12361 43004
rect 12065 42950 12111 43002
rect 12111 42950 12121 43002
rect 12145 42950 12175 43002
rect 12175 42950 12187 43002
rect 12187 42950 12201 43002
rect 12225 42950 12239 43002
rect 12239 42950 12251 43002
rect 12251 42950 12281 43002
rect 12305 42950 12315 43002
rect 12315 42950 12361 43002
rect 12065 42948 12121 42950
rect 12145 42948 12201 42950
rect 12225 42948 12281 42950
rect 12305 42948 12361 42950
rect 11978 42590 12034 42646
rect 12438 42318 12494 42374
rect 4291 41914 4347 41916
rect 4371 41914 4427 41916
rect 4451 41914 4507 41916
rect 4531 41914 4587 41916
rect 4291 41862 4337 41914
rect 4337 41862 4347 41914
rect 4371 41862 4401 41914
rect 4401 41862 4413 41914
rect 4413 41862 4427 41914
rect 4451 41862 4465 41914
rect 4465 41862 4477 41914
rect 4477 41862 4507 41914
rect 4531 41862 4541 41914
rect 4541 41862 4587 41914
rect 4291 41860 4347 41862
rect 4371 41860 4427 41862
rect 4451 41860 4507 41862
rect 4531 41860 4587 41862
rect 12065 41914 12121 41916
rect 12145 41914 12201 41916
rect 12225 41914 12281 41916
rect 12305 41914 12361 41916
rect 12065 41862 12111 41914
rect 12111 41862 12121 41914
rect 12145 41862 12175 41914
rect 12175 41862 12187 41914
rect 12187 41862 12201 41914
rect 12225 41862 12239 41914
rect 12239 41862 12251 41914
rect 12251 41862 12281 41914
rect 12305 41862 12315 41914
rect 12315 41862 12361 41914
rect 12065 41860 12121 41862
rect 12145 41860 12201 41862
rect 12225 41860 12281 41862
rect 12305 41860 12361 41862
rect 11886 41774 11942 41830
rect 2134 41094 2190 41150
rect 4342 41094 4398 41150
rect 8178 41370 8234 41372
rect 8258 41370 8314 41372
rect 8338 41370 8394 41372
rect 8418 41370 8474 41372
rect 8178 41318 8224 41370
rect 8224 41318 8234 41370
rect 8258 41318 8288 41370
rect 8288 41318 8300 41370
rect 8300 41318 8314 41370
rect 8338 41318 8352 41370
rect 8352 41318 8364 41370
rect 8364 41318 8394 41370
rect 8418 41318 8428 41370
rect 8428 41318 8474 41370
rect 8178 41316 8234 41318
rect 8258 41316 8314 41318
rect 8338 41316 8394 41318
rect 8418 41316 8474 41318
rect 11702 41230 11758 41286
rect 6550 41094 6606 41150
rect 8022 41094 8078 41150
rect 11794 41094 11850 41150
rect 212 40826 508 40828
rect 212 40774 508 40826
rect 212 40772 508 40774
rect 4291 40826 4347 40828
rect 4371 40826 4427 40828
rect 4451 40826 4507 40828
rect 4531 40826 4587 40828
rect 4291 40774 4337 40826
rect 4337 40774 4347 40826
rect 4371 40774 4401 40826
rect 4401 40774 4413 40826
rect 4413 40774 4427 40826
rect 4451 40774 4465 40826
rect 4465 40774 4477 40826
rect 4477 40774 4507 40826
rect 4531 40774 4541 40826
rect 4541 40774 4587 40826
rect 4291 40772 4347 40774
rect 4371 40772 4427 40774
rect 4451 40772 4507 40774
rect 4531 40772 4587 40774
rect 12065 40826 12121 40828
rect 12145 40826 12201 40828
rect 12225 40826 12281 40828
rect 12305 40826 12361 40828
rect 12065 40774 12111 40826
rect 12111 40774 12121 40826
rect 12145 40774 12175 40826
rect 12175 40774 12187 40826
rect 12187 40774 12201 40826
rect 12225 40774 12239 40826
rect 12239 40774 12251 40826
rect 12251 40774 12281 40826
rect 12305 40774 12315 40826
rect 12315 40774 12361 40826
rect 12065 40772 12121 40774
rect 12145 40772 12201 40774
rect 12225 40772 12281 40774
rect 12305 40772 12361 40774
rect 12990 42626 12992 42646
rect 12992 42626 13044 42646
rect 13044 42626 13046 42646
rect 12990 42590 13046 42626
rect 12530 41502 12586 41558
rect 13082 41658 13138 41694
rect 13082 41638 13084 41658
rect 13084 41638 13136 41658
rect 13136 41638 13138 41658
rect 13266 41638 13322 41694
rect 12990 41553 12992 41558
rect 12992 41553 13044 41558
rect 13044 41553 13046 41558
rect 12990 41502 13046 41553
rect 12622 41114 12678 41150
rect 12622 41094 12624 41114
rect 12624 41094 12676 41114
rect 12676 41094 12678 41114
rect 14002 43834 14058 43870
rect 14002 43814 14004 43834
rect 14004 43814 14056 43834
rect 14056 43814 14058 43834
rect 14186 43270 14242 43326
rect 14738 44358 14794 44414
rect 14370 42590 14426 42646
rect 14922 43290 14978 43326
rect 14922 43270 14924 43290
rect 14924 43270 14976 43290
rect 14976 43270 14978 43290
rect 14002 41538 14004 41558
rect 14004 41538 14056 41558
rect 14056 41538 14058 41558
rect 14002 41502 14058 41538
rect 14278 41130 14280 41150
rect 14280 41130 14332 41150
rect 14332 41130 14334 41150
rect 15750 42590 15806 42646
rect 15952 44634 16008 44636
rect 16032 44634 16088 44636
rect 16112 44634 16168 44636
rect 16192 44634 16248 44636
rect 15952 44582 15998 44634
rect 15998 44582 16008 44634
rect 16032 44582 16062 44634
rect 16062 44582 16074 44634
rect 16074 44582 16088 44634
rect 16112 44582 16126 44634
rect 16126 44582 16138 44634
rect 16138 44582 16168 44634
rect 16192 44582 16202 44634
rect 16202 44582 16248 44634
rect 15952 44580 16008 44582
rect 16032 44580 16088 44582
rect 16112 44580 16168 44582
rect 16192 44580 16248 44582
rect 25226 44766 25282 44822
rect 15952 43546 16008 43548
rect 16032 43546 16088 43548
rect 16112 43546 16168 43548
rect 16192 43546 16248 43548
rect 15952 43494 15998 43546
rect 15998 43494 16008 43546
rect 16032 43494 16062 43546
rect 16062 43494 16074 43546
rect 16074 43494 16088 43546
rect 16112 43494 16126 43546
rect 16126 43494 16138 43546
rect 16138 43494 16168 43546
rect 16192 43494 16202 43546
rect 16202 43494 16248 43546
rect 15952 43492 16008 43494
rect 16032 43492 16088 43494
rect 16112 43492 16168 43494
rect 16192 43492 16248 43494
rect 15952 42458 16008 42460
rect 16032 42458 16088 42460
rect 16112 42458 16168 42460
rect 16192 42458 16248 42460
rect 15952 42406 15998 42458
rect 15998 42406 16008 42458
rect 16032 42406 16062 42458
rect 16062 42406 16074 42458
rect 16074 42406 16088 42458
rect 16112 42406 16126 42458
rect 16126 42406 16138 42458
rect 16138 42406 16168 42458
rect 16192 42406 16202 42458
rect 16202 42406 16248 42458
rect 15952 42404 16008 42406
rect 16032 42404 16088 42406
rect 16112 42404 16168 42406
rect 16192 42404 16248 42406
rect 15106 41910 15162 41966
rect 15566 42082 15568 42102
rect 15568 42082 15620 42102
rect 15620 42082 15622 42102
rect 15198 41774 15254 41830
rect 14278 41094 14334 41130
rect 8178 40282 8234 40284
rect 8258 40282 8314 40284
rect 8338 40282 8394 40284
rect 8418 40282 8474 40284
rect 8178 40230 8224 40282
rect 8224 40230 8234 40282
rect 8258 40230 8288 40282
rect 8288 40230 8300 40282
rect 8300 40230 8314 40282
rect 8338 40230 8352 40282
rect 8352 40230 8364 40282
rect 8364 40230 8394 40282
rect 8418 40230 8428 40282
rect 8428 40230 8474 40282
rect 8178 40228 8234 40230
rect 8258 40228 8314 40230
rect 8338 40228 8394 40230
rect 8418 40228 8474 40230
rect 15566 42046 15622 42082
rect 15566 41094 15622 41150
rect 16210 42046 16266 42102
rect 17406 44358 17462 44414
rect 17130 43270 17186 43326
rect 17038 42726 17094 42782
rect 16486 41774 16542 41830
rect 15952 41370 16008 41372
rect 16032 41370 16088 41372
rect 16112 41370 16168 41372
rect 16192 41370 16248 41372
rect 15952 41318 15998 41370
rect 15998 41318 16008 41370
rect 16032 41318 16062 41370
rect 16062 41318 16074 41370
rect 16074 41318 16088 41370
rect 16112 41318 16126 41370
rect 16126 41318 16138 41370
rect 16138 41318 16168 41370
rect 16192 41318 16202 41370
rect 16202 41318 16248 41370
rect 15952 41316 16008 41318
rect 16032 41316 16088 41318
rect 16112 41316 16168 41318
rect 16192 41316 16248 41318
rect 16118 41094 16174 41150
rect 16854 41366 16910 41422
rect 17222 42182 17278 42238
rect 17130 42046 17186 42102
rect 17406 41910 17462 41966
rect 19839 44090 19895 44092
rect 19919 44090 19975 44092
rect 19999 44090 20055 44092
rect 20079 44090 20135 44092
rect 19839 44038 19885 44090
rect 19885 44038 19895 44090
rect 19919 44038 19949 44090
rect 19949 44038 19961 44090
rect 19961 44038 19975 44090
rect 19999 44038 20013 44090
rect 20013 44038 20025 44090
rect 20025 44038 20055 44090
rect 20079 44038 20089 44090
rect 20089 44038 20135 44090
rect 19839 44036 19895 44038
rect 19919 44036 19975 44038
rect 19999 44036 20055 44038
rect 20079 44036 20135 44038
rect 18234 42610 18290 42646
rect 18234 42590 18236 42610
rect 18236 42590 18288 42610
rect 18288 42590 18290 42610
rect 19430 42082 19432 42102
rect 19432 42082 19484 42102
rect 19484 42082 19486 42102
rect 19430 42046 19486 42082
rect 21730 43950 21786 44006
rect 19890 43134 19946 43190
rect 19839 43002 19895 43004
rect 19919 43002 19975 43004
rect 19999 43002 20055 43004
rect 20079 43002 20135 43004
rect 19839 42950 19885 43002
rect 19885 42950 19895 43002
rect 19919 42950 19949 43002
rect 19949 42950 19961 43002
rect 19961 42950 19975 43002
rect 19999 42950 20013 43002
rect 20013 42950 20025 43002
rect 20025 42950 20055 43002
rect 20079 42950 20089 43002
rect 20089 42950 20135 43002
rect 19839 42948 19895 42950
rect 19919 42948 19975 42950
rect 19999 42948 20055 42950
rect 20079 42948 20135 42950
rect 19798 42218 19800 42238
rect 19800 42218 19852 42238
rect 19852 42218 19854 42238
rect 19798 42182 19854 42218
rect 20258 42218 20260 42238
rect 20260 42218 20312 42238
rect 20312 42218 20314 42238
rect 20258 42182 20314 42218
rect 19839 41914 19895 41916
rect 19919 41914 19975 41916
rect 19999 41914 20055 41916
rect 20079 41914 20135 41916
rect 19839 41862 19885 41914
rect 19885 41862 19895 41914
rect 19919 41862 19949 41914
rect 19949 41862 19961 41914
rect 19961 41862 19975 41914
rect 19999 41862 20013 41914
rect 20013 41862 20025 41914
rect 20025 41862 20055 41914
rect 20079 41862 20089 41914
rect 20089 41862 20135 41914
rect 19839 41860 19895 41862
rect 19919 41860 19975 41862
rect 19999 41860 20055 41862
rect 20079 41860 20135 41862
rect 17498 41502 17554 41558
rect 17314 41366 17370 41422
rect 20994 42182 21050 42238
rect 20810 42082 20812 42102
rect 20812 42082 20864 42102
rect 20864 42082 20866 42102
rect 20810 42046 20866 42082
rect 20350 41638 20406 41694
rect 17682 41094 17738 41150
rect 17958 41094 18014 41150
rect 20626 41094 20682 41150
rect 22466 43134 22522 43190
rect 22650 42182 22706 42238
rect 23726 44634 23782 44636
rect 23806 44634 23862 44636
rect 23886 44634 23942 44636
rect 23966 44634 24022 44636
rect 23726 44582 23772 44634
rect 23772 44582 23782 44634
rect 23806 44582 23836 44634
rect 23836 44582 23848 44634
rect 23848 44582 23862 44634
rect 23886 44582 23900 44634
rect 23900 44582 23912 44634
rect 23912 44582 23942 44634
rect 23966 44582 23976 44634
rect 23976 44582 24022 44634
rect 23726 44580 23782 44582
rect 23806 44580 23862 44582
rect 23886 44580 23942 44582
rect 23966 44580 24022 44582
rect 25502 44630 25558 44686
rect 26790 44630 26846 44686
rect 28630 44630 28686 44686
rect 23662 43970 23718 44006
rect 23662 43950 23664 43970
rect 23664 43950 23716 43970
rect 23716 43950 23718 43970
rect 23726 43546 23782 43548
rect 23806 43546 23862 43548
rect 23886 43546 23942 43548
rect 23966 43546 24022 43548
rect 23726 43494 23772 43546
rect 23772 43494 23782 43546
rect 23806 43494 23836 43546
rect 23836 43494 23848 43546
rect 23848 43494 23862 43546
rect 23886 43494 23900 43546
rect 23900 43494 23912 43546
rect 23912 43494 23942 43546
rect 23966 43494 23976 43546
rect 23976 43494 24022 43546
rect 23726 43492 23782 43494
rect 23806 43492 23862 43494
rect 23886 43492 23942 43494
rect 23966 43492 24022 43494
rect 21454 41538 21456 41558
rect 21456 41538 21508 41558
rect 21508 41538 21510 41558
rect 23726 42458 23782 42460
rect 23806 42458 23862 42460
rect 23886 42458 23942 42460
rect 23966 42458 24022 42460
rect 23726 42406 23772 42458
rect 23772 42406 23782 42458
rect 23806 42406 23836 42458
rect 23836 42406 23848 42458
rect 23848 42406 23862 42458
rect 23886 42406 23900 42458
rect 23900 42406 23912 42458
rect 23912 42406 23942 42458
rect 23966 42406 23976 42458
rect 23976 42406 24022 42458
rect 23726 42404 23782 42406
rect 23806 42404 23862 42406
rect 23886 42404 23942 42406
rect 23966 42404 24022 42406
rect 31500 44634 31556 44636
rect 31580 44634 31636 44636
rect 31660 44634 31716 44636
rect 31740 44634 31796 44636
rect 31500 44582 31546 44634
rect 31546 44582 31556 44634
rect 31580 44582 31610 44634
rect 31610 44582 31622 44634
rect 31622 44582 31636 44634
rect 31660 44582 31674 44634
rect 31674 44582 31686 44634
rect 31686 44582 31716 44634
rect 31740 44582 31750 44634
rect 31750 44582 31796 44634
rect 31500 44580 31556 44582
rect 31580 44580 31636 44582
rect 31660 44580 31716 44582
rect 31740 44580 31796 44582
rect 27613 44090 27669 44092
rect 27693 44090 27749 44092
rect 27773 44090 27829 44092
rect 27853 44090 27909 44092
rect 27613 44038 27659 44090
rect 27659 44038 27669 44090
rect 27693 44038 27723 44090
rect 27723 44038 27735 44090
rect 27735 44038 27749 44090
rect 27773 44038 27787 44090
rect 27787 44038 27799 44090
rect 27799 44038 27829 44090
rect 27853 44038 27863 44090
rect 27863 44038 27909 44090
rect 27613 44036 27669 44038
rect 27693 44036 27749 44038
rect 27773 44036 27829 44038
rect 27853 44036 27909 44038
rect 28078 44086 28134 44142
rect 28814 43814 28870 43870
rect 25226 43134 25282 43190
rect 26054 43170 26056 43190
rect 26056 43170 26108 43190
rect 26108 43170 26110 43190
rect 26054 43134 26110 43170
rect 27613 43002 27669 43004
rect 27693 43002 27749 43004
rect 27773 43002 27829 43004
rect 27853 43002 27909 43004
rect 27613 42950 27659 43002
rect 27659 42950 27669 43002
rect 27693 42950 27723 43002
rect 27723 42950 27735 43002
rect 27735 42950 27749 43002
rect 27773 42950 27787 43002
rect 27787 42950 27799 43002
rect 27799 42950 27829 43002
rect 27853 42950 27863 43002
rect 27863 42950 27909 43002
rect 27613 42948 27669 42950
rect 27693 42948 27749 42950
rect 27773 42948 27829 42950
rect 27853 42948 27909 42950
rect 29550 44086 29606 44142
rect 30930 43950 30986 44006
rect 31500 43546 31556 43548
rect 31580 43546 31636 43548
rect 31660 43546 31716 43548
rect 31740 43546 31796 43548
rect 31500 43494 31546 43546
rect 31546 43494 31556 43546
rect 31580 43494 31610 43546
rect 31610 43494 31622 43546
rect 31622 43494 31636 43546
rect 31660 43494 31674 43546
rect 31674 43494 31686 43546
rect 31686 43494 31716 43546
rect 31740 43494 31750 43546
rect 31750 43494 31796 43546
rect 31500 43492 31556 43494
rect 31580 43492 31636 43494
rect 31660 43492 31716 43494
rect 31740 43492 31796 43494
rect 31500 42458 31556 42460
rect 31580 42458 31636 42460
rect 31660 42458 31716 42460
rect 31740 42458 31796 42460
rect 31500 42406 31546 42458
rect 31546 42406 31556 42458
rect 31580 42406 31610 42458
rect 31610 42406 31622 42458
rect 31622 42406 31636 42458
rect 31660 42406 31674 42458
rect 31674 42406 31686 42458
rect 31686 42406 31716 42458
rect 31740 42406 31750 42458
rect 31750 42406 31796 42458
rect 31500 42404 31556 42406
rect 31580 42404 31636 42406
rect 31660 42404 31716 42406
rect 31740 42404 31796 42406
rect 27613 41914 27669 41916
rect 27693 41914 27749 41916
rect 27773 41914 27829 41916
rect 27853 41914 27909 41916
rect 27613 41862 27659 41914
rect 27659 41862 27669 41914
rect 27693 41862 27723 41914
rect 27723 41862 27735 41914
rect 27735 41862 27749 41914
rect 27773 41862 27787 41914
rect 27787 41862 27799 41914
rect 27799 41862 27829 41914
rect 27853 41862 27863 41914
rect 27863 41862 27909 41914
rect 27613 41860 27669 41862
rect 27693 41860 27749 41862
rect 27773 41860 27829 41862
rect 27853 41860 27909 41862
rect 30746 41774 30802 41830
rect 21454 41502 21510 41538
rect 23726 41370 23782 41372
rect 23806 41370 23862 41372
rect 23886 41370 23942 41372
rect 23966 41370 24022 41372
rect 23726 41318 23772 41370
rect 23772 41318 23782 41370
rect 23806 41318 23836 41370
rect 23836 41318 23848 41370
rect 23848 41318 23862 41370
rect 23886 41318 23900 41370
rect 23900 41318 23912 41370
rect 23912 41318 23942 41370
rect 23966 41318 23976 41370
rect 23976 41318 24022 41370
rect 23726 41316 23782 41318
rect 23806 41316 23862 41318
rect 23886 41316 23942 41318
rect 23966 41316 24022 41318
rect 22834 41130 22836 41150
rect 22836 41130 22888 41150
rect 22888 41130 22890 41150
rect 22834 41094 22890 41130
rect 23570 41114 23626 41150
rect 23570 41094 23572 41114
rect 23572 41094 23624 41114
rect 23624 41094 23626 41114
rect 25778 41094 25834 41150
rect 30194 41130 30196 41150
rect 30196 41130 30248 41150
rect 30248 41130 30250 41150
rect 31500 41370 31556 41372
rect 31580 41370 31636 41372
rect 31660 41370 31716 41372
rect 31740 41370 31796 41372
rect 31500 41318 31546 41370
rect 31546 41318 31556 41370
rect 31580 41318 31610 41370
rect 31610 41318 31622 41370
rect 31622 41318 31636 41370
rect 31660 41318 31674 41370
rect 31674 41318 31686 41370
rect 31686 41318 31716 41370
rect 31740 41318 31750 41370
rect 31750 41318 31796 41370
rect 31500 41316 31556 41318
rect 31580 41316 31636 41318
rect 31660 41316 31716 41318
rect 31740 41316 31796 41318
rect 30194 41094 30250 41130
rect 19839 40826 19895 40828
rect 19919 40826 19975 40828
rect 19999 40826 20055 40828
rect 20079 40826 20135 40828
rect 19839 40774 19885 40826
rect 19885 40774 19895 40826
rect 19919 40774 19949 40826
rect 19949 40774 19961 40826
rect 19961 40774 19975 40826
rect 19999 40774 20013 40826
rect 20013 40774 20025 40826
rect 20025 40774 20055 40826
rect 20079 40774 20089 40826
rect 20089 40774 20135 40826
rect 19839 40772 19895 40774
rect 19919 40772 19975 40774
rect 19999 40772 20055 40774
rect 20079 40772 20135 40774
rect 15952 40282 16008 40284
rect 16032 40282 16088 40284
rect 16112 40282 16168 40284
rect 16192 40282 16248 40284
rect 15952 40230 15998 40282
rect 15998 40230 16008 40282
rect 16032 40230 16062 40282
rect 16062 40230 16074 40282
rect 16074 40230 16088 40282
rect 16112 40230 16126 40282
rect 16126 40230 16138 40282
rect 16138 40230 16168 40282
rect 16192 40230 16202 40282
rect 16202 40230 16248 40282
rect 15952 40228 16008 40230
rect 16032 40228 16088 40230
rect 16112 40228 16168 40230
rect 16192 40228 16248 40230
rect 14370 40142 14426 40198
rect 27613 40826 27669 40828
rect 27693 40826 27749 40828
rect 27773 40826 27829 40828
rect 27853 40826 27909 40828
rect 27613 40774 27659 40826
rect 27659 40774 27669 40826
rect 27693 40774 27723 40826
rect 27723 40774 27735 40826
rect 27735 40774 27749 40826
rect 27773 40774 27787 40826
rect 27787 40774 27799 40826
rect 27799 40774 27829 40826
rect 27853 40774 27863 40826
rect 27863 40774 27909 40826
rect 27613 40772 27669 40774
rect 27693 40772 27749 40774
rect 27773 40772 27829 40774
rect 27853 40772 27909 40774
rect 23726 40282 23782 40284
rect 23806 40282 23862 40284
rect 23886 40282 23942 40284
rect 23966 40282 24022 40284
rect 23726 40230 23772 40282
rect 23772 40230 23782 40282
rect 23806 40230 23836 40282
rect 23836 40230 23848 40282
rect 23848 40230 23862 40282
rect 23886 40230 23900 40282
rect 23900 40230 23912 40282
rect 23912 40230 23942 40282
rect 23966 40230 23976 40282
rect 23976 40230 24022 40282
rect 27250 40278 27306 40334
rect 23726 40228 23782 40230
rect 23806 40228 23862 40230
rect 23886 40228 23942 40230
rect 23966 40228 24022 40230
rect 31500 40282 31556 40284
rect 31580 40282 31636 40284
rect 31660 40282 31716 40284
rect 31740 40282 31796 40284
rect 31500 40230 31546 40282
rect 31546 40230 31556 40282
rect 31580 40230 31610 40282
rect 31610 40230 31622 40282
rect 31622 40230 31636 40282
rect 31660 40230 31674 40282
rect 31674 40230 31686 40282
rect 31686 40230 31716 40282
rect 31740 40230 31750 40282
rect 31750 40230 31796 40282
rect 31500 40228 31556 40230
rect 31580 40228 31636 40230
rect 31660 40228 31716 40230
rect 31740 40228 31796 40230
rect 28722 40142 28778 40198
rect 8148 39968 8502 40048
rect 12806 40006 12862 40062
rect 16946 40006 17002 40062
rect 1058 39740 1150 39792
rect 1058 39736 1150 39740
rect 2980 39736 3072 39792
rect 542 39606 598 39662
rect 31410 39606 31466 39662
rect 607 39474 663 39530
rect 31345 39474 31401 39530
rect 672 39342 728 39398
rect 31280 39342 31336 39398
rect 737 39210 793 39266
rect 31215 39210 31271 39266
rect 802 39078 858 39134
rect 31150 39078 31206 39134
rect 867 38946 923 39002
rect 31085 38946 31141 39002
rect 932 38814 988 38870
rect 31020 38814 31076 38870
rect 997 38682 1053 38738
rect 30955 38682 31011 38738
rect 1062 38550 1118 38606
rect 30890 38550 30946 38606
rect 1127 38418 1183 38474
rect 30825 38418 30881 38474
rect 1192 38286 1248 38342
rect 30760 38286 30816 38342
rect 1257 38154 1313 38210
rect 30695 38154 30751 38210
rect 1322 38022 1378 38078
rect 30630 38022 30686 38078
rect 1387 37890 1443 37946
rect 30565 37890 30621 37946
rect 1452 37758 1508 37814
rect 30500 37758 30556 37814
rect 1517 37626 1573 37682
rect 30435 37626 30491 37682
rect 1582 37494 1638 37550
rect 30370 37494 30426 37550
rect 5073 31496 5265 31688
rect 26732 31495 26924 31687
rect 5073 29496 5265 29688
rect 26732 29495 26924 29687
rect 31546 39494 31760 39752
rect 31760 39494 31764 39752
rect 5073 27496 5265 27688
rect 26732 27495 26924 27687
rect 5073 25496 5265 25688
rect 26732 25495 26924 25687
rect 5073 23496 5265 23688
rect 26732 23495 26924 23687
rect 5073 21496 5265 21688
rect 26732 21495 26924 21687
rect 5073 19496 5265 19688
rect 26732 19495 26924 19687
rect 5073 17496 5265 17688
rect 26732 17495 26924 17687
rect 5073 15496 5265 15688
rect 26732 15495 26924 15687
rect 5073 13496 5265 13688
rect 26732 13495 26924 13687
rect 5073 11496 5265 11688
rect 26732 11495 26924 11687
rect 5073 9496 5265 9688
rect 26732 9495 26924 9687
rect 5073 7496 5265 7688
rect 26732 7495 26924 7687
rect 5073 5496 5265 5688
rect 26732 5495 26924 5687
rect 5073 3496 5265 3688
rect 26732 3495 26924 3687
rect 5073 1496 5265 1688
rect 26732 1495 26924 1687
<< metal3 >>
rect 4521 44826 4587 44827
rect 4470 44762 4476 44826
rect 4540 44824 4587 44826
rect 15837 44824 15903 44827
rect 16246 44824 16252 44826
rect 4540 44822 4632 44824
rect 4582 44766 4632 44822
rect 4540 44764 4632 44766
rect 15837 44822 16252 44824
rect 15837 44766 15842 44822
rect 15898 44766 16252 44822
rect 15837 44764 16252 44766
rect 4540 44762 4587 44764
rect 4521 44761 4587 44762
rect 15837 44761 15903 44764
rect 16246 44762 16252 44764
rect 16316 44762 16322 44826
rect 17033 44824 17099 44827
rect 17718 44824 17724 44826
rect 17033 44822 17724 44824
rect 17033 44766 17038 44822
rect 17094 44766 17724 44822
rect 17033 44764 17724 44766
rect 17033 44761 17099 44764
rect 17718 44762 17724 44764
rect 17788 44762 17794 44826
rect 24342 44762 24348 44826
rect 24412 44824 24418 44826
rect 25221 44824 25287 44827
rect 24412 44822 25287 44824
rect 24412 44766 25226 44822
rect 25282 44766 25287 44822
rect 24412 44764 25287 44766
rect 24412 44762 24418 44764
rect 25221 44761 25287 44764
rect 9673 44690 9739 44691
rect 9622 44688 9628 44690
rect 8168 44640 8484 44641
rect 8168 44576 8174 44640
rect 8238 44576 8254 44640
rect 8318 44576 8334 44640
rect 8398 44576 8414 44640
rect 8478 44576 8484 44640
rect 9582 44628 9628 44688
rect 9692 44686 9739 44690
rect 9734 44630 9739 44686
rect 9622 44626 9628 44628
rect 9692 44626 9739 44630
rect 9673 44625 9739 44626
rect 15942 44640 16258 44641
rect 8168 44575 8484 44576
rect 15942 44576 15948 44640
rect 16012 44576 16028 44640
rect 16092 44576 16108 44640
rect 16172 44576 16188 44640
rect 16252 44576 16258 44640
rect 15942 44575 16258 44576
rect 23716 44640 24032 44641
rect 23716 44576 23722 44640
rect 23786 44576 23802 44640
rect 23866 44576 23882 44640
rect 23946 44576 23962 44640
rect 24026 44576 24032 44640
rect 25078 44626 25084 44690
rect 25148 44688 25154 44690
rect 25497 44688 25563 44691
rect 25148 44686 25563 44688
rect 25148 44630 25502 44686
rect 25558 44630 25563 44686
rect 25148 44628 25563 44630
rect 25148 44626 25154 44628
rect 25497 44625 25563 44628
rect 26550 44626 26556 44690
rect 26620 44688 26626 44690
rect 26785 44688 26851 44691
rect 26620 44686 26851 44688
rect 26620 44630 26790 44686
rect 26846 44630 26851 44686
rect 26620 44628 26851 44630
rect 26620 44626 26626 44628
rect 26785 44625 26851 44628
rect 27286 44626 27292 44690
rect 27356 44688 27362 44690
rect 28625 44688 28691 44691
rect 27356 44686 28691 44688
rect 27356 44630 28630 44686
rect 28686 44630 28691 44686
rect 27356 44628 28691 44630
rect 27356 44626 27362 44628
rect 28625 44625 28691 44628
rect 31490 44640 31806 44641
rect 23716 44575 24032 44576
rect 31490 44576 31496 44640
rect 31560 44576 31576 44640
rect 31640 44576 31656 44640
rect 31720 44576 31736 44640
rect 31800 44576 31806 44640
rect 31490 44575 31806 44576
rect 841 44554 907 44555
rect 1577 44554 1643 44555
rect 2313 44554 2379 44555
rect 790 44490 796 44554
rect 860 44552 907 44554
rect 860 44550 952 44552
rect 902 44494 952 44550
rect 860 44492 952 44494
rect 860 44490 907 44492
rect 1526 44490 1532 44554
rect 1596 44552 1643 44554
rect 1596 44550 1688 44552
rect 1638 44494 1688 44550
rect 1596 44492 1688 44494
rect 1596 44490 1643 44492
rect 2262 44490 2268 44554
rect 2332 44552 2379 44554
rect 2332 44550 2424 44552
rect 2374 44494 2424 44550
rect 2332 44492 2424 44494
rect 2332 44490 2379 44492
rect 2998 44490 3004 44554
rect 3068 44552 3074 44554
rect 3233 44552 3299 44555
rect 3785 44554 3851 44555
rect 5257 44554 5323 44555
rect 5993 44554 6059 44555
rect 3068 44550 3299 44552
rect 3068 44494 3238 44550
rect 3294 44494 3299 44550
rect 3068 44492 3299 44494
rect 3068 44490 3074 44492
rect 841 44489 907 44490
rect 1577 44489 1643 44490
rect 2313 44489 2379 44490
rect 3233 44489 3299 44492
rect 3734 44490 3740 44554
rect 3804 44552 3851 44554
rect 3804 44550 3896 44552
rect 3846 44494 3896 44550
rect 3804 44492 3896 44494
rect 3804 44490 3851 44492
rect 5206 44490 5212 44554
rect 5276 44552 5323 44554
rect 5276 44550 5368 44552
rect 5318 44494 5368 44550
rect 5276 44492 5368 44494
rect 5276 44490 5323 44492
rect 5942 44490 5948 44554
rect 6012 44552 6059 44554
rect 6012 44550 6104 44552
rect 6054 44494 6104 44550
rect 6012 44492 6104 44494
rect 6012 44490 6059 44492
rect 12566 44490 12572 44554
rect 12636 44552 12642 44554
rect 14089 44552 14155 44555
rect 12636 44550 14155 44552
rect 12636 44494 14094 44550
rect 14150 44494 14155 44550
rect 12636 44492 14155 44494
rect 12636 44490 12642 44492
rect 3785 44489 3851 44490
rect 5257 44489 5323 44490
rect 5993 44489 6059 44490
rect 14089 44489 14155 44492
rect 14733 44416 14799 44419
rect 15510 44416 15516 44418
rect 14733 44414 15516 44416
rect 14733 44358 14738 44414
rect 14794 44358 15516 44414
rect 14733 44356 15516 44358
rect 14733 44353 14799 44356
rect 15510 44354 15516 44356
rect 15580 44354 15586 44418
rect 16982 44354 16988 44418
rect 17052 44416 17058 44418
rect 17401 44416 17467 44419
rect 17052 44414 17467 44416
rect 17052 44358 17406 44414
rect 17462 44358 17467 44414
rect 17052 44356 17467 44358
rect 17052 44354 17058 44356
rect 17401 44353 17467 44356
rect 28073 44146 28139 44147
rect 29545 44146 29611 44147
rect 202 44096 518 44097
rect 202 44032 208 44096
rect 512 44032 518 44096
rect 202 44031 518 44032
rect 4281 44096 4597 44097
rect 4281 44032 4287 44096
rect 4351 44032 4367 44096
rect 4431 44032 4447 44096
rect 4511 44032 4527 44096
rect 4591 44032 4597 44096
rect 4281 44031 4597 44032
rect 12055 44096 12371 44097
rect 12055 44032 12061 44096
rect 12125 44032 12141 44096
rect 12205 44032 12221 44096
rect 12285 44032 12301 44096
rect 12365 44032 12371 44096
rect 12055 44031 12371 44032
rect 19829 44096 20145 44097
rect 19829 44032 19835 44096
rect 19899 44032 19915 44096
rect 19979 44032 19995 44096
rect 20059 44032 20075 44096
rect 20139 44032 20145 44096
rect 19829 44031 20145 44032
rect 27603 44096 27919 44097
rect 27603 44032 27609 44096
rect 27673 44032 27689 44096
rect 27753 44032 27769 44096
rect 27833 44032 27849 44096
rect 27913 44032 27919 44096
rect 28022 44082 28028 44146
rect 28092 44144 28139 44146
rect 29494 44144 29500 44146
rect 28092 44142 28184 44144
rect 28134 44086 28184 44142
rect 28092 44084 28184 44086
rect 29454 44084 29500 44144
rect 29564 44142 29611 44146
rect 29606 44086 29611 44142
rect 28092 44082 28139 44084
rect 29494 44082 29500 44084
rect 29564 44082 29611 44086
rect 28073 44081 28139 44082
rect 29545 44081 29611 44082
rect 27603 44031 27919 44032
rect 21725 44008 21791 44011
rect 23657 44008 23723 44011
rect 21725 44006 23723 44008
rect 21725 43950 21730 44006
rect 21786 43950 23662 44006
rect 23718 43950 23723 44006
rect 21725 43948 23723 43950
rect 21725 43945 21791 43948
rect 23657 43945 23723 43948
rect 30925 44010 30991 44011
rect 30925 44006 30972 44010
rect 31036 44008 31042 44010
rect 30925 43950 30930 44006
rect 30925 43946 30972 43950
rect 31036 43948 31082 44008
rect 31036 43946 31042 43948
rect 30925 43945 30991 43946
rect 13997 43874 14063 43875
rect 28809 43874 28875 43875
rect 13997 43872 14044 43874
rect 13952 43870 14044 43872
rect 13952 43814 14002 43870
rect 13952 43812 14044 43814
rect 13997 43810 14044 43812
rect 14108 43810 14114 43874
rect 28758 43872 28764 43874
rect 28718 43812 28764 43872
rect 28828 43870 28875 43874
rect 28870 43814 28875 43870
rect 28758 43810 28764 43812
rect 28828 43810 28875 43814
rect 13997 43809 14063 43810
rect 28809 43809 28875 43810
rect 8168 43552 8484 43553
rect 8168 43488 8174 43552
rect 8238 43488 8254 43552
rect 8318 43488 8334 43552
rect 8398 43488 8414 43552
rect 8478 43488 8484 43552
rect 8168 43487 8484 43488
rect 15942 43552 16258 43553
rect 15942 43488 15948 43552
rect 16012 43488 16028 43552
rect 16092 43488 16108 43552
rect 16172 43488 16188 43552
rect 16252 43488 16258 43552
rect 15942 43487 16258 43488
rect 23716 43552 24032 43553
rect 23716 43488 23722 43552
rect 23786 43488 23802 43552
rect 23866 43488 23882 43552
rect 23946 43488 23962 43552
rect 24026 43488 24032 43552
rect 23716 43487 24032 43488
rect 31490 43552 31806 43553
rect 31490 43488 31496 43552
rect 31560 43488 31576 43552
rect 31640 43488 31656 43552
rect 31720 43488 31736 43552
rect 31800 43488 31806 43552
rect 31490 43487 31806 43488
rect 14181 43328 14247 43331
rect 14774 43328 14780 43330
rect 14181 43326 14780 43328
rect 14181 43270 14186 43326
rect 14242 43270 14780 43326
rect 14181 43268 14780 43270
rect 14181 43265 14247 43268
rect 14774 43266 14780 43268
rect 14844 43266 14850 43330
rect 14917 43328 14983 43331
rect 17125 43328 17191 43331
rect 14917 43326 17191 43328
rect 14917 43270 14922 43326
rect 14978 43270 17130 43326
rect 17186 43270 17191 43326
rect 14917 43268 17191 43270
rect 14917 43265 14983 43268
rect 17125 43265 17191 43268
rect 19885 43192 19951 43195
rect 22461 43192 22527 43195
rect 25221 43192 25287 43195
rect 26049 43192 26115 43195
rect 19885 43190 26115 43192
rect 19885 43134 19890 43190
rect 19946 43134 22466 43190
rect 22522 43134 25226 43190
rect 25282 43134 26054 43190
rect 26110 43134 26115 43190
rect 19885 43132 26115 43134
rect 19885 43129 19951 43132
rect 22461 43129 22527 43132
rect 25221 43129 25287 43132
rect 26049 43129 26115 43132
rect 202 43008 518 43009
rect 202 42944 208 43008
rect 512 42944 518 43008
rect 202 42943 518 42944
rect 4281 43008 4597 43009
rect 4281 42944 4287 43008
rect 4351 42944 4367 43008
rect 4431 42944 4447 43008
rect 4511 42944 4527 43008
rect 4591 42944 4597 43008
rect 4281 42943 4597 42944
rect 12055 43008 12371 43009
rect 12055 42944 12061 43008
rect 12125 42944 12141 43008
rect 12205 42944 12221 43008
rect 12285 42944 12301 43008
rect 12365 42944 12371 43008
rect 12055 42943 12371 42944
rect 19829 43008 20145 43009
rect 19829 42944 19835 43008
rect 19899 42944 19915 43008
rect 19979 42944 19995 43008
rect 20059 42944 20075 43008
rect 20139 42944 20145 43008
rect 19829 42943 20145 42944
rect 27603 43008 27919 43009
rect 27603 42944 27609 43008
rect 27673 42944 27689 43008
rect 27753 42944 27769 43008
rect 27833 42944 27849 43008
rect 27913 42944 27919 43008
rect 27603 42943 27919 42944
rect 11145 42784 11211 42787
rect 17033 42784 17099 42787
rect 11145 42782 17099 42784
rect 11145 42726 11150 42782
rect 11206 42726 17038 42782
rect 17094 42726 17099 42782
rect 11145 42724 17099 42726
rect 11145 42721 11211 42724
rect 17033 42721 17099 42724
rect 11973 42648 12039 42651
rect 12985 42648 13051 42651
rect 11973 42646 13051 42648
rect 11973 42590 11978 42646
rect 12034 42590 12990 42646
rect 13046 42590 13051 42646
rect 11973 42588 13051 42590
rect 11973 42585 12039 42588
rect 12985 42585 13051 42588
rect 14365 42648 14431 42651
rect 15745 42648 15811 42651
rect 18229 42648 18295 42651
rect 14365 42646 18295 42648
rect 14365 42590 14370 42646
rect 14426 42590 15750 42646
rect 15806 42590 18234 42646
rect 18290 42590 18295 42646
rect 14365 42588 18295 42590
rect 14365 42585 14431 42588
rect 15745 42585 15811 42588
rect 18229 42585 18295 42588
rect 8168 42464 8484 42465
rect 8168 42400 8174 42464
rect 8238 42400 8254 42464
rect 8318 42400 8334 42464
rect 8398 42400 8414 42464
rect 8478 42400 8484 42464
rect 8168 42399 8484 42400
rect 15942 42464 16258 42465
rect 15942 42400 15948 42464
rect 16012 42400 16028 42464
rect 16092 42400 16108 42464
rect 16172 42400 16188 42464
rect 16252 42400 16258 42464
rect 15942 42399 16258 42400
rect 23716 42464 24032 42465
rect 23716 42400 23722 42464
rect 23786 42400 23802 42464
rect 23866 42400 23882 42464
rect 23946 42400 23962 42464
rect 24026 42400 24032 42464
rect 23716 42399 24032 42400
rect 31490 42464 31806 42465
rect 31490 42400 31496 42464
rect 31560 42400 31576 42464
rect 31640 42400 31656 42464
rect 31720 42400 31736 42464
rect 31800 42400 31806 42464
rect 31490 42399 31806 42400
rect 12433 42376 12499 42379
rect 13302 42376 13308 42378
rect 12433 42374 13308 42376
rect 12433 42318 12438 42374
rect 12494 42318 13308 42374
rect 12433 42316 13308 42318
rect 12433 42313 12499 42316
rect 13302 42314 13308 42316
rect 13372 42314 13378 42378
rect 7414 42178 7420 42242
rect 7484 42240 7490 42242
rect 11145 42240 11211 42243
rect 17217 42240 17283 42243
rect 7484 42238 11211 42240
rect 7484 42182 11150 42238
rect 11206 42182 11211 42238
rect 7484 42180 11211 42182
rect 7484 42178 7490 42180
rect 11145 42177 11211 42180
rect 11286 42238 17283 42240
rect 11286 42182 17222 42238
rect 17278 42182 17283 42238
rect 11286 42180 17283 42182
rect 11286 42107 11346 42180
rect 17217 42177 17283 42180
rect 19793 42240 19859 42243
rect 20253 42240 20319 42243
rect 20989 42240 21055 42243
rect 19793 42238 21055 42240
rect 19793 42182 19798 42238
rect 19854 42182 20258 42238
rect 20314 42182 20994 42238
rect 21050 42182 21055 42238
rect 19793 42180 21055 42182
rect 19793 42177 19859 42180
rect 20253 42177 20319 42180
rect 20989 42177 21055 42180
rect 22645 42240 22711 42243
rect 30230 42240 30236 42242
rect 22645 42238 30236 42240
rect 22645 42182 22650 42238
rect 22706 42182 30236 42238
rect 22645 42180 30236 42182
rect 22645 42177 22711 42180
rect 30230 42178 30236 42180
rect 30300 42178 30306 42242
rect 7966 42042 7972 42106
rect 8036 42104 8042 42106
rect 11237 42104 11346 42107
rect 15561 42104 15627 42107
rect 8036 42102 11346 42104
rect 8036 42046 11242 42102
rect 11298 42046 11346 42102
rect 8036 42044 11346 42046
rect 11470 42102 15627 42104
rect 11470 42046 15566 42102
rect 15622 42046 15627 42102
rect 11470 42044 15627 42046
rect 8036 42042 8042 42044
rect 11237 42041 11303 42044
rect 202 41920 518 41921
rect 202 41856 208 41920
rect 512 41856 518 41920
rect 202 41855 518 41856
rect 4281 41920 4597 41921
rect 4281 41856 4287 41920
rect 4351 41856 4367 41920
rect 4431 41856 4447 41920
rect 4511 41856 4527 41920
rect 4591 41856 4597 41920
rect 10358 41906 10364 41970
rect 10428 41968 10434 41970
rect 11470 41968 11530 42044
rect 15561 42041 15627 42044
rect 16205 42104 16271 42107
rect 17125 42104 17191 42107
rect 16205 42102 17191 42104
rect 16205 42046 16210 42102
rect 16266 42046 17130 42102
rect 17186 42046 17191 42102
rect 16205 42044 17191 42046
rect 16205 42041 16271 42044
rect 17125 42041 17191 42044
rect 19425 42104 19491 42107
rect 20805 42104 20871 42107
rect 19425 42102 20871 42104
rect 19425 42046 19430 42102
rect 19486 42046 20810 42102
rect 20866 42046 20871 42102
rect 19425 42044 20871 42046
rect 19425 42041 19491 42044
rect 20805 42041 20871 42044
rect 10428 41908 11530 41968
rect 15101 41968 15167 41971
rect 17401 41968 17467 41971
rect 15101 41966 17467 41968
rect 12055 41920 12371 41921
rect 10428 41906 10434 41908
rect 4281 41855 4597 41856
rect 12055 41856 12061 41920
rect 12125 41856 12141 41920
rect 12205 41856 12221 41920
rect 12285 41856 12301 41920
rect 12365 41856 12371 41920
rect 15101 41910 15106 41966
rect 15162 41910 17406 41966
rect 17462 41910 17467 41966
rect 15101 41908 17467 41910
rect 15101 41905 15167 41908
rect 17401 41905 17467 41908
rect 19829 41920 20145 41921
rect 12055 41855 12371 41856
rect 19829 41856 19835 41920
rect 19899 41856 19915 41920
rect 19979 41856 19995 41920
rect 20059 41856 20075 41920
rect 20139 41856 20145 41920
rect 19829 41855 20145 41856
rect 27603 41920 27919 41921
rect 27603 41856 27609 41920
rect 27673 41856 27689 41920
rect 27753 41856 27769 41920
rect 27833 41856 27849 41920
rect 27913 41856 27919 41920
rect 27603 41855 27919 41856
rect 8886 41770 8892 41834
rect 8956 41832 8962 41834
rect 11881 41832 11947 41835
rect 8956 41830 11947 41832
rect 8956 41774 11886 41830
rect 11942 41774 11947 41830
rect 8956 41772 11947 41774
rect 8956 41770 8962 41772
rect 11881 41769 11947 41772
rect 15193 41832 15259 41835
rect 16481 41832 16547 41835
rect 15193 41830 16547 41832
rect 15193 41774 15198 41830
rect 15254 41774 16486 41830
rect 16542 41774 16547 41830
rect 15193 41772 16547 41774
rect 15193 41769 15259 41772
rect 16481 41769 16547 41772
rect 30741 41832 30807 41835
rect 31334 41832 31340 41834
rect 30741 41830 31340 41832
rect 30741 41774 30746 41830
rect 30802 41774 31340 41830
rect 30741 41772 31340 41774
rect 30741 41769 30807 41772
rect 31334 41770 31340 41772
rect 31404 41770 31410 41834
rect 6678 41634 6684 41698
rect 6748 41696 6754 41698
rect 13077 41696 13143 41699
rect 6748 41694 13143 41696
rect 6748 41638 13082 41694
rect 13138 41638 13143 41694
rect 6748 41636 13143 41638
rect 6748 41634 6754 41636
rect 13077 41633 13143 41636
rect 13261 41696 13327 41699
rect 20345 41696 20411 41699
rect 13261 41694 20411 41696
rect 13261 41638 13266 41694
rect 13322 41638 20350 41694
rect 20406 41638 20411 41694
rect 13261 41636 20411 41638
rect 13261 41633 13327 41636
rect 20345 41633 20411 41636
rect 4654 41498 4660 41562
rect 4724 41560 4730 41562
rect 12525 41560 12591 41563
rect 4724 41558 12591 41560
rect 4724 41502 12530 41558
rect 12586 41502 12591 41558
rect 4724 41500 12591 41502
rect 4724 41498 4730 41500
rect 12525 41497 12591 41500
rect 12985 41560 13051 41563
rect 13997 41560 14063 41563
rect 17493 41560 17559 41563
rect 21449 41560 21515 41563
rect 12985 41558 14063 41560
rect 12985 41502 12990 41558
rect 13046 41502 14002 41558
rect 14058 41502 14063 41558
rect 12985 41500 14063 41502
rect 12985 41497 13051 41500
rect 13997 41497 14063 41500
rect 15748 41558 21515 41560
rect 15748 41502 17498 41558
rect 17554 41502 21454 41558
rect 21510 41502 21515 41558
rect 15748 41500 21515 41502
rect 8168 41376 8484 41377
rect 8168 41312 8174 41376
rect 8238 41312 8254 41376
rect 8318 41312 8334 41376
rect 8398 41312 8414 41376
rect 8478 41312 8484 41376
rect 11094 41362 11100 41426
rect 11164 41424 11170 41426
rect 15748 41424 15808 41500
rect 17493 41497 17559 41500
rect 21449 41497 21515 41500
rect 11164 41364 15808 41424
rect 16849 41424 16915 41427
rect 17309 41424 17375 41427
rect 16849 41422 17375 41424
rect 15942 41376 16258 41377
rect 11164 41362 11170 41364
rect 8168 41311 8484 41312
rect 15942 41312 15948 41376
rect 16012 41312 16028 41376
rect 16092 41312 16108 41376
rect 16172 41312 16188 41376
rect 16252 41312 16258 41376
rect 16849 41366 16854 41422
rect 16910 41366 17314 41422
rect 17370 41366 17375 41422
rect 16849 41364 17375 41366
rect 16849 41361 16915 41364
rect 17309 41361 17375 41364
rect 23716 41376 24032 41377
rect 15942 41311 16258 41312
rect 23716 41312 23722 41376
rect 23786 41312 23802 41376
rect 23866 41312 23882 41376
rect 23946 41312 23962 41376
rect 24026 41312 24032 41376
rect 23716 41311 24032 41312
rect 31490 41376 31806 41377
rect 31490 41312 31496 41376
rect 31560 41312 31576 41376
rect 31640 41312 31656 41376
rect 31720 41312 31736 41376
rect 31800 41312 31806 41376
rect 31490 41311 31806 41312
rect 9622 41226 9628 41290
rect 9692 41288 9698 41290
rect 11697 41288 11763 41291
rect 9692 41286 11763 41288
rect 9692 41230 11702 41286
rect 11758 41230 11763 41286
rect 9692 41228 11763 41230
rect 9692 41226 9698 41228
rect 11697 41225 11763 41228
rect 11830 41226 11836 41290
rect 11900 41288 11906 41290
rect 11900 41228 15808 41288
rect 11900 41226 11906 41228
rect 1342 41090 1348 41154
rect 1412 41152 1418 41154
rect 2129 41152 2195 41155
rect 1412 41150 2195 41152
rect 1412 41094 2134 41150
rect 2190 41094 2195 41150
rect 1412 41092 2195 41094
rect 1412 41090 1418 41092
rect 2129 41089 2195 41092
rect 2814 41090 2820 41154
rect 2884 41152 2890 41154
rect 4337 41152 4403 41155
rect 2884 41150 4403 41152
rect 2884 41094 4342 41150
rect 4398 41094 4403 41150
rect 2884 41092 4403 41094
rect 2884 41090 2890 41092
rect 4337 41089 4403 41092
rect 5758 41090 5764 41154
rect 5828 41152 5834 41154
rect 6545 41152 6611 41155
rect 5828 41150 6611 41152
rect 5828 41094 6550 41150
rect 6606 41094 6611 41150
rect 5828 41092 6611 41094
rect 5828 41090 5834 41092
rect 6545 41089 6611 41092
rect 7230 41090 7236 41154
rect 7300 41152 7306 41154
rect 8017 41152 8083 41155
rect 7300 41150 8083 41152
rect 7300 41094 8022 41150
rect 8078 41094 8083 41150
rect 7300 41092 8083 41094
rect 7300 41090 7306 41092
rect 8017 41089 8083 41092
rect 11094 41090 11100 41154
rect 11164 41152 11170 41154
rect 11789 41152 11855 41155
rect 11164 41150 11855 41152
rect 11164 41094 11794 41150
rect 11850 41094 11855 41150
rect 11164 41092 11855 41094
rect 11164 41090 11170 41092
rect 11789 41089 11855 41092
rect 12617 41152 12683 41155
rect 14273 41152 14339 41155
rect 15561 41154 15627 41155
rect 15510 41152 15516 41154
rect 12617 41150 14339 41152
rect 12617 41094 12622 41150
rect 12678 41094 14278 41150
rect 14334 41094 14339 41150
rect 12617 41092 14339 41094
rect 15470 41092 15516 41152
rect 15580 41150 15627 41154
rect 15622 41094 15627 41150
rect 12617 41089 12683 41092
rect 14273 41089 14339 41092
rect 15510 41090 15516 41092
rect 15580 41090 15627 41094
rect 15748 41152 15808 41228
rect 16113 41152 16179 41155
rect 17677 41152 17743 41155
rect 15748 41150 17743 41152
rect 15748 41094 16118 41150
rect 16174 41094 17682 41150
rect 17738 41094 17743 41150
rect 15748 41092 17743 41094
rect 15561 41089 15627 41090
rect 16113 41089 16179 41092
rect 17677 41089 17743 41092
rect 17953 41152 18019 41155
rect 18454 41152 18460 41154
rect 17953 41150 18460 41152
rect 17953 41094 17958 41150
rect 18014 41094 18460 41150
rect 17953 41092 18460 41094
rect 17953 41089 18019 41092
rect 18454 41090 18460 41092
rect 18524 41090 18530 41154
rect 20621 41152 20687 41155
rect 22829 41154 22895 41155
rect 21398 41152 21404 41154
rect 20621 41150 21404 41152
rect 20621 41094 20626 41150
rect 20682 41094 21404 41150
rect 20621 41092 21404 41094
rect 20621 41089 20687 41092
rect 21398 41090 21404 41092
rect 21468 41090 21474 41154
rect 22829 41150 22876 41154
rect 22940 41152 22946 41154
rect 23565 41152 23631 41155
rect 25773 41154 25839 41155
rect 30189 41154 30255 41155
rect 24342 41152 24348 41154
rect 22829 41094 22834 41150
rect 22829 41090 22876 41094
rect 22940 41092 22986 41152
rect 23565 41150 24348 41152
rect 23565 41094 23570 41150
rect 23626 41094 24348 41150
rect 23565 41092 24348 41094
rect 22940 41090 22946 41092
rect 22829 41089 22895 41090
rect 23565 41089 23631 41092
rect 24342 41090 24348 41092
rect 24412 41090 24418 41154
rect 25773 41150 25820 41154
rect 25884 41152 25890 41154
rect 25773 41094 25778 41150
rect 25773 41090 25820 41094
rect 25884 41092 25930 41152
rect 30189 41150 30236 41154
rect 30300 41152 30306 41154
rect 30189 41094 30194 41150
rect 25884 41090 25890 41092
rect 30189 41090 30236 41094
rect 30300 41092 30346 41152
rect 30300 41090 30306 41092
rect 25773 41089 25839 41090
rect 30189 41089 30255 41090
rect 202 40832 518 40833
rect 202 40768 208 40832
rect 512 40768 518 40832
rect 202 40767 518 40768
rect 4281 40832 4597 40833
rect 4281 40768 4287 40832
rect 4351 40768 4367 40832
rect 4431 40768 4447 40832
rect 4511 40768 4527 40832
rect 4591 40768 4597 40832
rect 4281 40767 4597 40768
rect 12055 40832 12371 40833
rect 12055 40768 12061 40832
rect 12125 40768 12141 40832
rect 12205 40768 12221 40832
rect 12285 40768 12301 40832
rect 12365 40768 12371 40832
rect 12055 40767 12371 40768
rect 19829 40832 20145 40833
rect 19829 40768 19835 40832
rect 19899 40768 19915 40832
rect 19979 40768 19995 40832
rect 20059 40768 20075 40832
rect 20139 40768 20145 40832
rect 19829 40767 20145 40768
rect 27603 40832 27919 40833
rect 27603 40768 27609 40832
rect 27673 40768 27689 40832
rect 27753 40768 27769 40832
rect 27833 40768 27849 40832
rect 27913 40768 27919 40832
rect 27603 40767 27919 40768
rect 27245 40338 27311 40339
rect 27245 40334 27292 40338
rect 27356 40336 27362 40338
rect 8168 40288 8484 40289
rect 8168 40224 8174 40288
rect 8238 40224 8254 40288
rect 8318 40224 8334 40288
rect 8398 40224 8414 40288
rect 8478 40224 8484 40288
rect 8168 40223 8484 40224
rect 15942 40288 16258 40289
rect 15942 40224 15948 40288
rect 16012 40224 16028 40288
rect 16092 40224 16108 40288
rect 16172 40224 16188 40288
rect 16252 40224 16258 40288
rect 15942 40223 16258 40224
rect 23716 40288 24032 40289
rect 23716 40224 23722 40288
rect 23786 40224 23802 40288
rect 23866 40224 23882 40288
rect 23946 40224 23962 40288
rect 24026 40224 24032 40288
rect 27245 40278 27250 40334
rect 27245 40274 27292 40278
rect 27356 40276 27402 40336
rect 31490 40288 31806 40289
rect 27356 40274 27362 40276
rect 27245 40273 27311 40274
rect 23716 40223 24032 40224
rect 31490 40224 31496 40288
rect 31560 40224 31576 40288
rect 31640 40224 31656 40288
rect 31720 40224 31736 40288
rect 31800 40224 31806 40288
rect 31490 40223 31806 40224
rect 14038 40138 14044 40202
rect 14108 40200 14114 40202
rect 14365 40200 14431 40203
rect 14108 40198 14431 40200
rect 14108 40142 14370 40198
rect 14426 40142 14431 40198
rect 14108 40140 14431 40142
rect 14108 40138 14114 40140
rect 14365 40137 14431 40140
rect 28717 40202 28783 40203
rect 28717 40198 28764 40202
rect 28828 40200 28834 40202
rect 28717 40142 28722 40198
rect 28717 40138 28764 40142
rect 28828 40140 28874 40200
rect 28828 40138 28834 40140
rect 28717 40137 28783 40138
rect 8128 40048 8178 40054
rect 8472 40048 8522 40054
rect 8128 39968 8148 40048
rect 8502 39968 8522 40048
rect 12566 40002 12572 40066
rect 12636 40064 12642 40066
rect 12801 40064 12867 40067
rect 12636 40062 12867 40064
rect 12636 40006 12806 40062
rect 12862 40006 12867 40062
rect 12636 40004 12867 40006
rect 12636 40002 12642 40004
rect 12801 40001 12867 40004
rect 16941 40066 17007 40067
rect 16941 40062 16988 40066
rect 17052 40064 17058 40066
rect 16941 40006 16946 40062
rect 16941 40002 16988 40006
rect 17052 40004 17098 40064
rect 17052 40002 17058 40004
rect 16941 40001 17007 40002
rect 8128 39962 8178 39968
rect 8472 39962 8522 39968
rect 1050 39796 1158 39802
rect 1376 39796 1454 39803
rect 1050 39792 1454 39796
rect 1050 39736 1058 39792
rect 1150 39736 1454 39792
rect 1050 39726 1158 39736
rect 1376 39725 1454 39736
rect 2848 39802 2926 39804
rect 2848 39798 3080 39802
rect 2848 39731 2854 39798
rect 2920 39792 3080 39798
rect 2920 39736 2980 39792
rect 3072 39736 3080 39792
rect 2920 39731 3080 39736
rect 2848 39726 3080 39731
rect 31534 39758 31776 39764
rect 2848 39725 2926 39726
rect 30229 39670 30305 39674
rect 534 39664 606 39670
rect 30229 39664 30235 39670
rect 534 39662 30235 39664
rect 534 39606 542 39662
rect 598 39606 30235 39662
rect 30299 39664 30305 39670
rect 31402 39664 31474 39670
rect 30299 39662 31474 39664
rect 30299 39606 31410 39662
rect 31466 39606 31474 39662
rect 534 39604 31474 39606
rect 534 39598 606 39604
rect 31402 39598 31474 39604
rect 28757 39538 28833 39542
rect 599 39532 671 39538
rect 28757 39532 28763 39538
rect 599 39530 28763 39532
rect 599 39474 607 39530
rect 663 39474 28763 39530
rect 28827 39532 28833 39538
rect 31337 39532 31409 39538
rect 28827 39530 31410 39532
rect 28827 39474 31345 39530
rect 31401 39474 31410 39530
rect 31534 39488 31540 39758
rect 31770 39488 31776 39758
rect 31534 39482 31776 39488
rect 599 39472 31410 39474
rect 599 39466 671 39472
rect 31337 39466 31409 39472
rect 27285 39406 27361 39410
rect 664 39400 736 39406
rect 27285 39400 27291 39406
rect 664 39398 27291 39400
rect 664 39342 672 39398
rect 728 39342 27291 39398
rect 27355 39400 27361 39406
rect 31272 39400 31344 39406
rect 27355 39398 31345 39400
rect 27355 39342 31280 39398
rect 31336 39342 31345 39398
rect 664 39340 31345 39342
rect 664 39334 736 39340
rect 31272 39334 31344 39340
rect 25813 39274 25889 39278
rect 729 39268 801 39274
rect 25813 39268 25819 39274
rect 729 39266 25819 39268
rect 729 39210 737 39266
rect 793 39210 25819 39266
rect 25883 39268 25889 39274
rect 31207 39268 31279 39274
rect 25883 39266 31280 39268
rect 25883 39210 31215 39266
rect 31271 39210 31280 39266
rect 729 39208 31280 39210
rect 729 39202 801 39208
rect 31207 39202 31279 39208
rect 24341 39142 24417 39146
rect 794 39136 866 39142
rect 24341 39136 24347 39142
rect 794 39134 24347 39136
rect 794 39078 802 39134
rect 858 39078 24347 39134
rect 24411 39136 24417 39142
rect 31142 39136 31214 39142
rect 24411 39134 31215 39136
rect 24411 39078 31150 39134
rect 31206 39078 31215 39134
rect 794 39076 31215 39078
rect 794 39070 866 39076
rect 31142 39070 31214 39076
rect 22869 39010 22945 39014
rect 859 39004 931 39010
rect 22869 39004 22875 39010
rect 859 39002 22875 39004
rect 859 38946 867 39002
rect 923 38946 22875 39002
rect 22939 39004 22945 39010
rect 31077 39004 31149 39010
rect 22939 39002 31150 39004
rect 22939 38946 31085 39002
rect 31141 38946 31150 39002
rect 859 38944 31150 38946
rect 859 38938 931 38944
rect 31077 38938 31149 38944
rect 21397 38878 21473 38882
rect 924 38872 996 38878
rect 21397 38872 21403 38878
rect 924 38870 21403 38872
rect 924 38814 932 38870
rect 988 38814 21403 38870
rect 21467 38872 21473 38878
rect 31012 38872 31084 38878
rect 21467 38870 31085 38872
rect 21467 38814 31020 38870
rect 31076 38814 31085 38870
rect 924 38812 31085 38814
rect 924 38806 996 38812
rect 31012 38806 31084 38812
rect 18453 38746 18529 38750
rect 989 38740 1061 38746
rect 18453 38740 18459 38746
rect 989 38738 18459 38740
rect 989 38682 997 38738
rect 1053 38682 18459 38738
rect 18523 38740 18529 38746
rect 30947 38740 31019 38746
rect 18523 38738 31020 38740
rect 18523 38682 30955 38738
rect 31011 38682 31020 38738
rect 989 38680 31020 38682
rect 989 38674 1061 38680
rect 30947 38674 31019 38680
rect 16981 38614 17057 38618
rect 1054 38608 1126 38614
rect 16981 38608 16987 38614
rect 1054 38606 16987 38608
rect 1054 38550 1062 38606
rect 1118 38550 16987 38606
rect 17051 38608 17057 38614
rect 30882 38608 30954 38614
rect 17051 38606 30955 38608
rect 17051 38550 30890 38606
rect 30946 38550 30955 38606
rect 1054 38548 30955 38550
rect 1054 38542 1126 38548
rect 30882 38542 30954 38548
rect 15509 38482 15585 38486
rect 1119 38476 1191 38482
rect 15509 38476 15515 38482
rect 1119 38474 15515 38476
rect 1119 38418 1127 38474
rect 1183 38418 15515 38474
rect 15579 38476 15585 38482
rect 30817 38476 30889 38482
rect 15579 38474 30890 38476
rect 15579 38418 30825 38474
rect 30881 38418 30890 38474
rect 1119 38416 30890 38418
rect 1119 38410 1191 38416
rect 30817 38410 30889 38416
rect 14037 38350 14113 38354
rect 1184 38344 1256 38350
rect 14037 38344 14043 38350
rect 1184 38342 14043 38344
rect 1184 38286 1192 38342
rect 1248 38286 14043 38342
rect 14107 38344 14113 38350
rect 30752 38344 30824 38350
rect 14107 38342 30825 38344
rect 14107 38286 30760 38342
rect 30816 38286 30825 38342
rect 1184 38284 30825 38286
rect 1184 38278 1256 38284
rect 30752 38278 30824 38284
rect 12565 38218 12641 38222
rect 1249 38212 1321 38218
rect 12565 38212 12571 38218
rect 1249 38210 12571 38212
rect 1249 38154 1257 38210
rect 1313 38154 12571 38210
rect 12635 38212 12641 38218
rect 30687 38212 30759 38218
rect 12635 38210 30760 38212
rect 12635 38154 30695 38210
rect 30751 38154 30760 38210
rect 1249 38152 30760 38154
rect 1249 38146 1321 38152
rect 30687 38146 30759 38152
rect 11093 38086 11169 38090
rect 1314 38080 1386 38086
rect 11093 38080 11099 38086
rect 1314 38078 11099 38080
rect 1314 38022 1322 38078
rect 1378 38022 11099 38078
rect 11163 38080 11169 38086
rect 30622 38080 30694 38086
rect 11163 38078 30695 38080
rect 11163 38022 30630 38078
rect 30686 38022 30695 38078
rect 1314 38020 30695 38022
rect 1314 38014 1386 38020
rect 30622 38014 30694 38020
rect 9621 37954 9697 37958
rect 1379 37948 1451 37954
rect 9621 37948 9627 37954
rect 1379 37946 9627 37948
rect 1379 37890 1387 37946
rect 1443 37890 9627 37946
rect 9691 37948 9697 37954
rect 30557 37948 30629 37954
rect 9691 37946 30630 37948
rect 9691 37890 30565 37946
rect 30621 37890 30630 37946
rect 1379 37888 30630 37890
rect 1379 37882 1451 37888
rect 30557 37882 30629 37888
rect 7265 37822 7341 37826
rect 1444 37816 1516 37822
rect 7265 37816 7271 37822
rect 1444 37814 7271 37816
rect 1444 37758 1452 37814
rect 1508 37758 7271 37814
rect 7335 37816 7341 37822
rect 30492 37816 30564 37822
rect 7335 37814 30565 37816
rect 7335 37758 30500 37814
rect 30556 37758 30565 37814
rect 1444 37756 30565 37758
rect 1444 37750 1516 37756
rect 30492 37750 30564 37756
rect 5793 37690 5869 37694
rect 1509 37684 1581 37690
rect 5793 37684 5799 37690
rect 1509 37682 5799 37684
rect 1509 37626 1517 37682
rect 1573 37626 5799 37682
rect 5863 37684 5869 37690
rect 30427 37684 30499 37690
rect 5863 37682 30500 37684
rect 5863 37626 30435 37682
rect 30491 37626 30500 37682
rect 1509 37624 30500 37626
rect 1509 37618 1581 37624
rect 30427 37618 30499 37624
rect 4321 37558 4397 37562
rect 1574 37552 1646 37558
rect 4321 37552 4327 37558
rect 1574 37550 4327 37552
rect 1574 37494 1582 37550
rect 1638 37494 4327 37550
rect 4391 37552 4397 37558
rect 30362 37552 30434 37558
rect 4391 37550 30435 37552
rect 4391 37494 30370 37550
rect 30426 37494 30435 37550
rect 1574 37492 30435 37494
rect 1574 37486 1646 37492
rect 30362 37486 30434 37492
rect 5066 31689 5272 31695
rect 5066 31495 5072 31689
rect 5266 31495 5272 31689
rect 5066 31489 5272 31495
rect 26725 31688 26931 31694
rect 26725 31494 26731 31688
rect 26925 31494 26931 31688
rect 26725 31488 26931 31494
rect 5066 29689 5272 29695
rect 5066 29495 5072 29689
rect 5266 29495 5272 29689
rect 5066 29489 5272 29495
rect 26725 29688 26931 29694
rect 26725 29494 26731 29688
rect 26925 29494 26931 29688
rect 26725 29488 26931 29494
rect 5066 27689 5272 27695
rect 5066 27495 5072 27689
rect 5266 27495 5272 27689
rect 5066 27489 5272 27495
rect 26725 27688 26931 27694
rect 26725 27494 26731 27688
rect 26925 27494 26931 27688
rect 26725 27488 26931 27494
rect 5066 25689 5272 25695
rect 5066 25495 5072 25689
rect 5266 25495 5272 25689
rect 5066 25489 5272 25495
rect 26725 25688 26931 25694
rect 26725 25494 26731 25688
rect 26925 25494 26931 25688
rect 26725 25488 26931 25494
rect 5066 23689 5272 23695
rect 5066 23495 5072 23689
rect 5266 23495 5272 23689
rect 5066 23489 5272 23495
rect 26725 23688 26931 23694
rect 26725 23494 26731 23688
rect 26925 23494 26931 23688
rect 26725 23488 26931 23494
rect 5066 21689 5272 21695
rect 5066 21495 5072 21689
rect 5266 21495 5272 21689
rect 5066 21489 5272 21495
rect 26725 21688 26931 21694
rect 26725 21494 26731 21688
rect 26925 21494 26931 21688
rect 26725 21488 26931 21494
rect 5066 19689 5272 19695
rect 5066 19495 5072 19689
rect 5266 19495 5272 19689
rect 5066 19489 5272 19495
rect 26725 19688 26931 19694
rect 26725 19494 26731 19688
rect 26925 19494 26931 19688
rect 26725 19488 26931 19494
rect 5066 17689 5272 17695
rect 5066 17495 5072 17689
rect 5266 17495 5272 17689
rect 5066 17489 5272 17495
rect 26725 17688 26931 17694
rect 26725 17494 26731 17688
rect 26925 17494 26931 17688
rect 26725 17488 26931 17494
rect 5066 15689 5272 15695
rect 5066 15495 5072 15689
rect 5266 15495 5272 15689
rect 5066 15489 5272 15495
rect 26725 15688 26931 15694
rect 26725 15494 26731 15688
rect 26925 15494 26931 15688
rect 26725 15488 26931 15494
rect 5066 13689 5272 13695
rect 5066 13495 5072 13689
rect 5266 13495 5272 13689
rect 5066 13489 5272 13495
rect 26725 13688 26931 13694
rect 26725 13494 26731 13688
rect 26925 13494 26931 13688
rect 26725 13488 26931 13494
rect 5066 11689 5272 11695
rect 5066 11495 5072 11689
rect 5266 11495 5272 11689
rect 5066 11489 5272 11495
rect 26725 11688 26931 11694
rect 26725 11494 26731 11688
rect 26925 11494 26931 11688
rect 26725 11488 26931 11494
rect 5066 9689 5272 9695
rect 5066 9495 5072 9689
rect 5266 9495 5272 9689
rect 5066 9489 5272 9495
rect 26725 9688 26931 9694
rect 26725 9494 26731 9688
rect 26925 9494 26931 9688
rect 26725 9488 26931 9494
rect 5066 7689 5272 7695
rect 5066 7495 5072 7689
rect 5266 7495 5272 7689
rect 5066 7489 5272 7495
rect 26725 7688 26931 7694
rect 26725 7494 26731 7688
rect 26925 7494 26931 7688
rect 26725 7488 26931 7494
rect 5066 5689 5272 5695
rect 5066 5495 5072 5689
rect 5266 5495 5272 5689
rect 5066 5489 5272 5495
rect 26725 5688 26931 5694
rect 26725 5494 26731 5688
rect 26925 5494 26931 5688
rect 26725 5488 26931 5494
rect 5066 3689 5272 3695
rect 5066 3495 5072 3689
rect 5266 3495 5272 3689
rect 5066 3489 5272 3495
rect 26725 3688 26931 3694
rect 26725 3494 26731 3688
rect 26925 3494 26931 3688
rect 26725 3488 26931 3494
rect 5066 1689 5272 1695
rect 5066 1495 5072 1689
rect 5266 1495 5272 1689
rect 5066 1489 5272 1495
rect 26725 1688 26931 1694
rect 26725 1494 26731 1688
rect 26925 1494 26931 1688
rect 26725 1488 26931 1494
<< via3 >>
rect 4476 44822 4540 44826
rect 4476 44766 4526 44822
rect 4526 44766 4540 44822
rect 4476 44762 4540 44766
rect 16252 44762 16316 44826
rect 17724 44762 17788 44826
rect 24348 44762 24412 44826
rect 8174 44636 8238 44640
rect 8174 44580 8178 44636
rect 8178 44580 8234 44636
rect 8234 44580 8238 44636
rect 8174 44576 8238 44580
rect 8254 44636 8318 44640
rect 8254 44580 8258 44636
rect 8258 44580 8314 44636
rect 8314 44580 8318 44636
rect 8254 44576 8318 44580
rect 8334 44636 8398 44640
rect 8334 44580 8338 44636
rect 8338 44580 8394 44636
rect 8394 44580 8398 44636
rect 8334 44576 8398 44580
rect 8414 44636 8478 44640
rect 8414 44580 8418 44636
rect 8418 44580 8474 44636
rect 8474 44580 8478 44636
rect 8414 44576 8478 44580
rect 9628 44686 9692 44690
rect 9628 44630 9678 44686
rect 9678 44630 9692 44686
rect 9628 44626 9692 44630
rect 15948 44636 16012 44640
rect 15948 44580 15952 44636
rect 15952 44580 16008 44636
rect 16008 44580 16012 44636
rect 15948 44576 16012 44580
rect 16028 44636 16092 44640
rect 16028 44580 16032 44636
rect 16032 44580 16088 44636
rect 16088 44580 16092 44636
rect 16028 44576 16092 44580
rect 16108 44636 16172 44640
rect 16108 44580 16112 44636
rect 16112 44580 16168 44636
rect 16168 44580 16172 44636
rect 16108 44576 16172 44580
rect 16188 44636 16252 44640
rect 16188 44580 16192 44636
rect 16192 44580 16248 44636
rect 16248 44580 16252 44636
rect 16188 44576 16252 44580
rect 23722 44636 23786 44640
rect 23722 44580 23726 44636
rect 23726 44580 23782 44636
rect 23782 44580 23786 44636
rect 23722 44576 23786 44580
rect 23802 44636 23866 44640
rect 23802 44580 23806 44636
rect 23806 44580 23862 44636
rect 23862 44580 23866 44636
rect 23802 44576 23866 44580
rect 23882 44636 23946 44640
rect 23882 44580 23886 44636
rect 23886 44580 23942 44636
rect 23942 44580 23946 44636
rect 23882 44576 23946 44580
rect 23962 44636 24026 44640
rect 23962 44580 23966 44636
rect 23966 44580 24022 44636
rect 24022 44580 24026 44636
rect 23962 44576 24026 44580
rect 25084 44626 25148 44690
rect 26556 44626 26620 44690
rect 27292 44626 27356 44690
rect 31496 44636 31560 44640
rect 31496 44580 31500 44636
rect 31500 44580 31556 44636
rect 31556 44580 31560 44636
rect 31496 44576 31560 44580
rect 31576 44636 31640 44640
rect 31576 44580 31580 44636
rect 31580 44580 31636 44636
rect 31636 44580 31640 44636
rect 31576 44576 31640 44580
rect 31656 44636 31720 44640
rect 31656 44580 31660 44636
rect 31660 44580 31716 44636
rect 31716 44580 31720 44636
rect 31656 44576 31720 44580
rect 31736 44636 31800 44640
rect 31736 44580 31740 44636
rect 31740 44580 31796 44636
rect 31796 44580 31800 44636
rect 31736 44576 31800 44580
rect 796 44550 860 44554
rect 796 44494 846 44550
rect 846 44494 860 44550
rect 796 44490 860 44494
rect 1532 44550 1596 44554
rect 1532 44494 1582 44550
rect 1582 44494 1596 44550
rect 1532 44490 1596 44494
rect 2268 44550 2332 44554
rect 2268 44494 2318 44550
rect 2318 44494 2332 44550
rect 2268 44490 2332 44494
rect 3004 44490 3068 44554
rect 3740 44550 3804 44554
rect 3740 44494 3790 44550
rect 3790 44494 3804 44550
rect 3740 44490 3804 44494
rect 5212 44550 5276 44554
rect 5212 44494 5262 44550
rect 5262 44494 5276 44550
rect 5212 44490 5276 44494
rect 5948 44550 6012 44554
rect 5948 44494 5998 44550
rect 5998 44494 6012 44550
rect 5948 44490 6012 44494
rect 12572 44490 12636 44554
rect 15516 44354 15580 44418
rect 16988 44354 17052 44418
rect 208 44092 512 44096
rect 208 44036 212 44092
rect 212 44036 508 44092
rect 508 44036 512 44092
rect 208 44032 512 44036
rect 4287 44092 4351 44096
rect 4287 44036 4291 44092
rect 4291 44036 4347 44092
rect 4347 44036 4351 44092
rect 4287 44032 4351 44036
rect 4367 44092 4431 44096
rect 4367 44036 4371 44092
rect 4371 44036 4427 44092
rect 4427 44036 4431 44092
rect 4367 44032 4431 44036
rect 4447 44092 4511 44096
rect 4447 44036 4451 44092
rect 4451 44036 4507 44092
rect 4507 44036 4511 44092
rect 4447 44032 4511 44036
rect 4527 44092 4591 44096
rect 4527 44036 4531 44092
rect 4531 44036 4587 44092
rect 4587 44036 4591 44092
rect 4527 44032 4591 44036
rect 12061 44092 12125 44096
rect 12061 44036 12065 44092
rect 12065 44036 12121 44092
rect 12121 44036 12125 44092
rect 12061 44032 12125 44036
rect 12141 44092 12205 44096
rect 12141 44036 12145 44092
rect 12145 44036 12201 44092
rect 12201 44036 12205 44092
rect 12141 44032 12205 44036
rect 12221 44092 12285 44096
rect 12221 44036 12225 44092
rect 12225 44036 12281 44092
rect 12281 44036 12285 44092
rect 12221 44032 12285 44036
rect 12301 44092 12365 44096
rect 12301 44036 12305 44092
rect 12305 44036 12361 44092
rect 12361 44036 12365 44092
rect 12301 44032 12365 44036
rect 19835 44092 19899 44096
rect 19835 44036 19839 44092
rect 19839 44036 19895 44092
rect 19895 44036 19899 44092
rect 19835 44032 19899 44036
rect 19915 44092 19979 44096
rect 19915 44036 19919 44092
rect 19919 44036 19975 44092
rect 19975 44036 19979 44092
rect 19915 44032 19979 44036
rect 19995 44092 20059 44096
rect 19995 44036 19999 44092
rect 19999 44036 20055 44092
rect 20055 44036 20059 44092
rect 19995 44032 20059 44036
rect 20075 44092 20139 44096
rect 20075 44036 20079 44092
rect 20079 44036 20135 44092
rect 20135 44036 20139 44092
rect 20075 44032 20139 44036
rect 27609 44092 27673 44096
rect 27609 44036 27613 44092
rect 27613 44036 27669 44092
rect 27669 44036 27673 44092
rect 27609 44032 27673 44036
rect 27689 44092 27753 44096
rect 27689 44036 27693 44092
rect 27693 44036 27749 44092
rect 27749 44036 27753 44092
rect 27689 44032 27753 44036
rect 27769 44092 27833 44096
rect 27769 44036 27773 44092
rect 27773 44036 27829 44092
rect 27829 44036 27833 44092
rect 27769 44032 27833 44036
rect 27849 44092 27913 44096
rect 27849 44036 27853 44092
rect 27853 44036 27909 44092
rect 27909 44036 27913 44092
rect 27849 44032 27913 44036
rect 28028 44142 28092 44146
rect 28028 44086 28078 44142
rect 28078 44086 28092 44142
rect 28028 44082 28092 44086
rect 29500 44142 29564 44146
rect 29500 44086 29550 44142
rect 29550 44086 29564 44142
rect 29500 44082 29564 44086
rect 30972 44006 31036 44010
rect 30972 43950 30986 44006
rect 30986 43950 31036 44006
rect 30972 43946 31036 43950
rect 14044 43870 14108 43874
rect 14044 43814 14058 43870
rect 14058 43814 14108 43870
rect 14044 43810 14108 43814
rect 28764 43870 28828 43874
rect 28764 43814 28814 43870
rect 28814 43814 28828 43870
rect 28764 43810 28828 43814
rect 8174 43548 8238 43552
rect 8174 43492 8178 43548
rect 8178 43492 8234 43548
rect 8234 43492 8238 43548
rect 8174 43488 8238 43492
rect 8254 43548 8318 43552
rect 8254 43492 8258 43548
rect 8258 43492 8314 43548
rect 8314 43492 8318 43548
rect 8254 43488 8318 43492
rect 8334 43548 8398 43552
rect 8334 43492 8338 43548
rect 8338 43492 8394 43548
rect 8394 43492 8398 43548
rect 8334 43488 8398 43492
rect 8414 43548 8478 43552
rect 8414 43492 8418 43548
rect 8418 43492 8474 43548
rect 8474 43492 8478 43548
rect 8414 43488 8478 43492
rect 15948 43548 16012 43552
rect 15948 43492 15952 43548
rect 15952 43492 16008 43548
rect 16008 43492 16012 43548
rect 15948 43488 16012 43492
rect 16028 43548 16092 43552
rect 16028 43492 16032 43548
rect 16032 43492 16088 43548
rect 16088 43492 16092 43548
rect 16028 43488 16092 43492
rect 16108 43548 16172 43552
rect 16108 43492 16112 43548
rect 16112 43492 16168 43548
rect 16168 43492 16172 43548
rect 16108 43488 16172 43492
rect 16188 43548 16252 43552
rect 16188 43492 16192 43548
rect 16192 43492 16248 43548
rect 16248 43492 16252 43548
rect 16188 43488 16252 43492
rect 23722 43548 23786 43552
rect 23722 43492 23726 43548
rect 23726 43492 23782 43548
rect 23782 43492 23786 43548
rect 23722 43488 23786 43492
rect 23802 43548 23866 43552
rect 23802 43492 23806 43548
rect 23806 43492 23862 43548
rect 23862 43492 23866 43548
rect 23802 43488 23866 43492
rect 23882 43548 23946 43552
rect 23882 43492 23886 43548
rect 23886 43492 23942 43548
rect 23942 43492 23946 43548
rect 23882 43488 23946 43492
rect 23962 43548 24026 43552
rect 23962 43492 23966 43548
rect 23966 43492 24022 43548
rect 24022 43492 24026 43548
rect 23962 43488 24026 43492
rect 31496 43548 31560 43552
rect 31496 43492 31500 43548
rect 31500 43492 31556 43548
rect 31556 43492 31560 43548
rect 31496 43488 31560 43492
rect 31576 43548 31640 43552
rect 31576 43492 31580 43548
rect 31580 43492 31636 43548
rect 31636 43492 31640 43548
rect 31576 43488 31640 43492
rect 31656 43548 31720 43552
rect 31656 43492 31660 43548
rect 31660 43492 31716 43548
rect 31716 43492 31720 43548
rect 31656 43488 31720 43492
rect 31736 43548 31800 43552
rect 31736 43492 31740 43548
rect 31740 43492 31796 43548
rect 31796 43492 31800 43548
rect 31736 43488 31800 43492
rect 14780 43266 14844 43330
rect 208 43004 512 43008
rect 208 42948 212 43004
rect 212 42948 508 43004
rect 508 42948 512 43004
rect 208 42944 512 42948
rect 4287 43004 4351 43008
rect 4287 42948 4291 43004
rect 4291 42948 4347 43004
rect 4347 42948 4351 43004
rect 4287 42944 4351 42948
rect 4367 43004 4431 43008
rect 4367 42948 4371 43004
rect 4371 42948 4427 43004
rect 4427 42948 4431 43004
rect 4367 42944 4431 42948
rect 4447 43004 4511 43008
rect 4447 42948 4451 43004
rect 4451 42948 4507 43004
rect 4507 42948 4511 43004
rect 4447 42944 4511 42948
rect 4527 43004 4591 43008
rect 4527 42948 4531 43004
rect 4531 42948 4587 43004
rect 4587 42948 4591 43004
rect 4527 42944 4591 42948
rect 12061 43004 12125 43008
rect 12061 42948 12065 43004
rect 12065 42948 12121 43004
rect 12121 42948 12125 43004
rect 12061 42944 12125 42948
rect 12141 43004 12205 43008
rect 12141 42948 12145 43004
rect 12145 42948 12201 43004
rect 12201 42948 12205 43004
rect 12141 42944 12205 42948
rect 12221 43004 12285 43008
rect 12221 42948 12225 43004
rect 12225 42948 12281 43004
rect 12281 42948 12285 43004
rect 12221 42944 12285 42948
rect 12301 43004 12365 43008
rect 12301 42948 12305 43004
rect 12305 42948 12361 43004
rect 12361 42948 12365 43004
rect 12301 42944 12365 42948
rect 19835 43004 19899 43008
rect 19835 42948 19839 43004
rect 19839 42948 19895 43004
rect 19895 42948 19899 43004
rect 19835 42944 19899 42948
rect 19915 43004 19979 43008
rect 19915 42948 19919 43004
rect 19919 42948 19975 43004
rect 19975 42948 19979 43004
rect 19915 42944 19979 42948
rect 19995 43004 20059 43008
rect 19995 42948 19999 43004
rect 19999 42948 20055 43004
rect 20055 42948 20059 43004
rect 19995 42944 20059 42948
rect 20075 43004 20139 43008
rect 20075 42948 20079 43004
rect 20079 42948 20135 43004
rect 20135 42948 20139 43004
rect 20075 42944 20139 42948
rect 27609 43004 27673 43008
rect 27609 42948 27613 43004
rect 27613 42948 27669 43004
rect 27669 42948 27673 43004
rect 27609 42944 27673 42948
rect 27689 43004 27753 43008
rect 27689 42948 27693 43004
rect 27693 42948 27749 43004
rect 27749 42948 27753 43004
rect 27689 42944 27753 42948
rect 27769 43004 27833 43008
rect 27769 42948 27773 43004
rect 27773 42948 27829 43004
rect 27829 42948 27833 43004
rect 27769 42944 27833 42948
rect 27849 43004 27913 43008
rect 27849 42948 27853 43004
rect 27853 42948 27909 43004
rect 27909 42948 27913 43004
rect 27849 42944 27913 42948
rect 8174 42460 8238 42464
rect 8174 42404 8178 42460
rect 8178 42404 8234 42460
rect 8234 42404 8238 42460
rect 8174 42400 8238 42404
rect 8254 42460 8318 42464
rect 8254 42404 8258 42460
rect 8258 42404 8314 42460
rect 8314 42404 8318 42460
rect 8254 42400 8318 42404
rect 8334 42460 8398 42464
rect 8334 42404 8338 42460
rect 8338 42404 8394 42460
rect 8394 42404 8398 42460
rect 8334 42400 8398 42404
rect 8414 42460 8478 42464
rect 8414 42404 8418 42460
rect 8418 42404 8474 42460
rect 8474 42404 8478 42460
rect 8414 42400 8478 42404
rect 15948 42460 16012 42464
rect 15948 42404 15952 42460
rect 15952 42404 16008 42460
rect 16008 42404 16012 42460
rect 15948 42400 16012 42404
rect 16028 42460 16092 42464
rect 16028 42404 16032 42460
rect 16032 42404 16088 42460
rect 16088 42404 16092 42460
rect 16028 42400 16092 42404
rect 16108 42460 16172 42464
rect 16108 42404 16112 42460
rect 16112 42404 16168 42460
rect 16168 42404 16172 42460
rect 16108 42400 16172 42404
rect 16188 42460 16252 42464
rect 16188 42404 16192 42460
rect 16192 42404 16248 42460
rect 16248 42404 16252 42460
rect 16188 42400 16252 42404
rect 23722 42460 23786 42464
rect 23722 42404 23726 42460
rect 23726 42404 23782 42460
rect 23782 42404 23786 42460
rect 23722 42400 23786 42404
rect 23802 42460 23866 42464
rect 23802 42404 23806 42460
rect 23806 42404 23862 42460
rect 23862 42404 23866 42460
rect 23802 42400 23866 42404
rect 23882 42460 23946 42464
rect 23882 42404 23886 42460
rect 23886 42404 23942 42460
rect 23942 42404 23946 42460
rect 23882 42400 23946 42404
rect 23962 42460 24026 42464
rect 23962 42404 23966 42460
rect 23966 42404 24022 42460
rect 24022 42404 24026 42460
rect 23962 42400 24026 42404
rect 31496 42460 31560 42464
rect 31496 42404 31500 42460
rect 31500 42404 31556 42460
rect 31556 42404 31560 42460
rect 31496 42400 31560 42404
rect 31576 42460 31640 42464
rect 31576 42404 31580 42460
rect 31580 42404 31636 42460
rect 31636 42404 31640 42460
rect 31576 42400 31640 42404
rect 31656 42460 31720 42464
rect 31656 42404 31660 42460
rect 31660 42404 31716 42460
rect 31716 42404 31720 42460
rect 31656 42400 31720 42404
rect 31736 42460 31800 42464
rect 31736 42404 31740 42460
rect 31740 42404 31796 42460
rect 31796 42404 31800 42460
rect 31736 42400 31800 42404
rect 13308 42314 13372 42378
rect 7420 42178 7484 42242
rect 30236 42178 30300 42242
rect 7972 42042 8036 42106
rect 208 41916 512 41920
rect 208 41860 212 41916
rect 212 41860 508 41916
rect 508 41860 512 41916
rect 208 41856 512 41860
rect 4287 41916 4351 41920
rect 4287 41860 4291 41916
rect 4291 41860 4347 41916
rect 4347 41860 4351 41916
rect 4287 41856 4351 41860
rect 4367 41916 4431 41920
rect 4367 41860 4371 41916
rect 4371 41860 4427 41916
rect 4427 41860 4431 41916
rect 4367 41856 4431 41860
rect 4447 41916 4511 41920
rect 4447 41860 4451 41916
rect 4451 41860 4507 41916
rect 4507 41860 4511 41916
rect 4447 41856 4511 41860
rect 4527 41916 4591 41920
rect 4527 41860 4531 41916
rect 4531 41860 4587 41916
rect 4587 41860 4591 41916
rect 4527 41856 4591 41860
rect 10364 41906 10428 41970
rect 12061 41916 12125 41920
rect 12061 41860 12065 41916
rect 12065 41860 12121 41916
rect 12121 41860 12125 41916
rect 12061 41856 12125 41860
rect 12141 41916 12205 41920
rect 12141 41860 12145 41916
rect 12145 41860 12201 41916
rect 12201 41860 12205 41916
rect 12141 41856 12205 41860
rect 12221 41916 12285 41920
rect 12221 41860 12225 41916
rect 12225 41860 12281 41916
rect 12281 41860 12285 41916
rect 12221 41856 12285 41860
rect 12301 41916 12365 41920
rect 12301 41860 12305 41916
rect 12305 41860 12361 41916
rect 12361 41860 12365 41916
rect 12301 41856 12365 41860
rect 19835 41916 19899 41920
rect 19835 41860 19839 41916
rect 19839 41860 19895 41916
rect 19895 41860 19899 41916
rect 19835 41856 19899 41860
rect 19915 41916 19979 41920
rect 19915 41860 19919 41916
rect 19919 41860 19975 41916
rect 19975 41860 19979 41916
rect 19915 41856 19979 41860
rect 19995 41916 20059 41920
rect 19995 41860 19999 41916
rect 19999 41860 20055 41916
rect 20055 41860 20059 41916
rect 19995 41856 20059 41860
rect 20075 41916 20139 41920
rect 20075 41860 20079 41916
rect 20079 41860 20135 41916
rect 20135 41860 20139 41916
rect 20075 41856 20139 41860
rect 27609 41916 27673 41920
rect 27609 41860 27613 41916
rect 27613 41860 27669 41916
rect 27669 41860 27673 41916
rect 27609 41856 27673 41860
rect 27689 41916 27753 41920
rect 27689 41860 27693 41916
rect 27693 41860 27749 41916
rect 27749 41860 27753 41916
rect 27689 41856 27753 41860
rect 27769 41916 27833 41920
rect 27769 41860 27773 41916
rect 27773 41860 27829 41916
rect 27829 41860 27833 41916
rect 27769 41856 27833 41860
rect 27849 41916 27913 41920
rect 27849 41860 27853 41916
rect 27853 41860 27909 41916
rect 27909 41860 27913 41916
rect 27849 41856 27913 41860
rect 8892 41770 8956 41834
rect 31340 41770 31404 41834
rect 6684 41634 6748 41698
rect 4660 41498 4724 41562
rect 8174 41372 8238 41376
rect 8174 41316 8178 41372
rect 8178 41316 8234 41372
rect 8234 41316 8238 41372
rect 8174 41312 8238 41316
rect 8254 41372 8318 41376
rect 8254 41316 8258 41372
rect 8258 41316 8314 41372
rect 8314 41316 8318 41372
rect 8254 41312 8318 41316
rect 8334 41372 8398 41376
rect 8334 41316 8338 41372
rect 8338 41316 8394 41372
rect 8394 41316 8398 41372
rect 8334 41312 8398 41316
rect 8414 41372 8478 41376
rect 8414 41316 8418 41372
rect 8418 41316 8474 41372
rect 8474 41316 8478 41372
rect 8414 41312 8478 41316
rect 11100 41362 11164 41426
rect 15948 41372 16012 41376
rect 15948 41316 15952 41372
rect 15952 41316 16008 41372
rect 16008 41316 16012 41372
rect 15948 41312 16012 41316
rect 16028 41372 16092 41376
rect 16028 41316 16032 41372
rect 16032 41316 16088 41372
rect 16088 41316 16092 41372
rect 16028 41312 16092 41316
rect 16108 41372 16172 41376
rect 16108 41316 16112 41372
rect 16112 41316 16168 41372
rect 16168 41316 16172 41372
rect 16108 41312 16172 41316
rect 16188 41372 16252 41376
rect 16188 41316 16192 41372
rect 16192 41316 16248 41372
rect 16248 41316 16252 41372
rect 16188 41312 16252 41316
rect 23722 41372 23786 41376
rect 23722 41316 23726 41372
rect 23726 41316 23782 41372
rect 23782 41316 23786 41372
rect 23722 41312 23786 41316
rect 23802 41372 23866 41376
rect 23802 41316 23806 41372
rect 23806 41316 23862 41372
rect 23862 41316 23866 41372
rect 23802 41312 23866 41316
rect 23882 41372 23946 41376
rect 23882 41316 23886 41372
rect 23886 41316 23942 41372
rect 23942 41316 23946 41372
rect 23882 41312 23946 41316
rect 23962 41372 24026 41376
rect 23962 41316 23966 41372
rect 23966 41316 24022 41372
rect 24022 41316 24026 41372
rect 23962 41312 24026 41316
rect 31496 41372 31560 41376
rect 31496 41316 31500 41372
rect 31500 41316 31556 41372
rect 31556 41316 31560 41372
rect 31496 41312 31560 41316
rect 31576 41372 31640 41376
rect 31576 41316 31580 41372
rect 31580 41316 31636 41372
rect 31636 41316 31640 41372
rect 31576 41312 31640 41316
rect 31656 41372 31720 41376
rect 31656 41316 31660 41372
rect 31660 41316 31716 41372
rect 31716 41316 31720 41372
rect 31656 41312 31720 41316
rect 31736 41372 31800 41376
rect 31736 41316 31740 41372
rect 31740 41316 31796 41372
rect 31796 41316 31800 41372
rect 31736 41312 31800 41316
rect 9628 41226 9692 41290
rect 11836 41226 11900 41290
rect 1348 41090 1412 41154
rect 2820 41090 2884 41154
rect 5764 41090 5828 41154
rect 7236 41090 7300 41154
rect 11100 41090 11164 41154
rect 15516 41150 15580 41154
rect 15516 41094 15566 41150
rect 15566 41094 15580 41150
rect 15516 41090 15580 41094
rect 18460 41090 18524 41154
rect 21404 41090 21468 41154
rect 22876 41150 22940 41154
rect 22876 41094 22890 41150
rect 22890 41094 22940 41150
rect 22876 41090 22940 41094
rect 24348 41090 24412 41154
rect 25820 41150 25884 41154
rect 25820 41094 25834 41150
rect 25834 41094 25884 41150
rect 25820 41090 25884 41094
rect 30236 41150 30300 41154
rect 30236 41094 30250 41150
rect 30250 41094 30300 41150
rect 30236 41090 30300 41094
rect 208 40828 512 40832
rect 208 40772 212 40828
rect 212 40772 508 40828
rect 508 40772 512 40828
rect 208 40768 512 40772
rect 4287 40828 4351 40832
rect 4287 40772 4291 40828
rect 4291 40772 4347 40828
rect 4347 40772 4351 40828
rect 4287 40768 4351 40772
rect 4367 40828 4431 40832
rect 4367 40772 4371 40828
rect 4371 40772 4427 40828
rect 4427 40772 4431 40828
rect 4367 40768 4431 40772
rect 4447 40828 4511 40832
rect 4447 40772 4451 40828
rect 4451 40772 4507 40828
rect 4507 40772 4511 40828
rect 4447 40768 4511 40772
rect 4527 40828 4591 40832
rect 4527 40772 4531 40828
rect 4531 40772 4587 40828
rect 4587 40772 4591 40828
rect 4527 40768 4591 40772
rect 12061 40828 12125 40832
rect 12061 40772 12065 40828
rect 12065 40772 12121 40828
rect 12121 40772 12125 40828
rect 12061 40768 12125 40772
rect 12141 40828 12205 40832
rect 12141 40772 12145 40828
rect 12145 40772 12201 40828
rect 12201 40772 12205 40828
rect 12141 40768 12205 40772
rect 12221 40828 12285 40832
rect 12221 40772 12225 40828
rect 12225 40772 12281 40828
rect 12281 40772 12285 40828
rect 12221 40768 12285 40772
rect 12301 40828 12365 40832
rect 12301 40772 12305 40828
rect 12305 40772 12361 40828
rect 12361 40772 12365 40828
rect 12301 40768 12365 40772
rect 19835 40828 19899 40832
rect 19835 40772 19839 40828
rect 19839 40772 19895 40828
rect 19895 40772 19899 40828
rect 19835 40768 19899 40772
rect 19915 40828 19979 40832
rect 19915 40772 19919 40828
rect 19919 40772 19975 40828
rect 19975 40772 19979 40828
rect 19915 40768 19979 40772
rect 19995 40828 20059 40832
rect 19995 40772 19999 40828
rect 19999 40772 20055 40828
rect 20055 40772 20059 40828
rect 19995 40768 20059 40772
rect 20075 40828 20139 40832
rect 20075 40772 20079 40828
rect 20079 40772 20135 40828
rect 20135 40772 20139 40828
rect 20075 40768 20139 40772
rect 27609 40828 27673 40832
rect 27609 40772 27613 40828
rect 27613 40772 27669 40828
rect 27669 40772 27673 40828
rect 27609 40768 27673 40772
rect 27689 40828 27753 40832
rect 27689 40772 27693 40828
rect 27693 40772 27749 40828
rect 27749 40772 27753 40828
rect 27689 40768 27753 40772
rect 27769 40828 27833 40832
rect 27769 40772 27773 40828
rect 27773 40772 27829 40828
rect 27829 40772 27833 40828
rect 27769 40768 27833 40772
rect 27849 40828 27913 40832
rect 27849 40772 27853 40828
rect 27853 40772 27909 40828
rect 27909 40772 27913 40828
rect 27849 40768 27913 40772
rect 27292 40334 27356 40338
rect 8174 40284 8238 40288
rect 8174 40228 8178 40284
rect 8178 40228 8234 40284
rect 8234 40228 8238 40284
rect 8174 40224 8238 40228
rect 8254 40284 8318 40288
rect 8254 40228 8258 40284
rect 8258 40228 8314 40284
rect 8314 40228 8318 40284
rect 8254 40224 8318 40228
rect 8334 40284 8398 40288
rect 8334 40228 8338 40284
rect 8338 40228 8394 40284
rect 8394 40228 8398 40284
rect 8334 40224 8398 40228
rect 8414 40284 8478 40288
rect 8414 40228 8418 40284
rect 8418 40228 8474 40284
rect 8474 40228 8478 40284
rect 8414 40224 8478 40228
rect 15948 40284 16012 40288
rect 15948 40228 15952 40284
rect 15952 40228 16008 40284
rect 16008 40228 16012 40284
rect 15948 40224 16012 40228
rect 16028 40284 16092 40288
rect 16028 40228 16032 40284
rect 16032 40228 16088 40284
rect 16088 40228 16092 40284
rect 16028 40224 16092 40228
rect 16108 40284 16172 40288
rect 16108 40228 16112 40284
rect 16112 40228 16168 40284
rect 16168 40228 16172 40284
rect 16108 40224 16172 40228
rect 16188 40284 16252 40288
rect 16188 40228 16192 40284
rect 16192 40228 16248 40284
rect 16248 40228 16252 40284
rect 16188 40224 16252 40228
rect 23722 40284 23786 40288
rect 23722 40228 23726 40284
rect 23726 40228 23782 40284
rect 23782 40228 23786 40284
rect 23722 40224 23786 40228
rect 23802 40284 23866 40288
rect 23802 40228 23806 40284
rect 23806 40228 23862 40284
rect 23862 40228 23866 40284
rect 23802 40224 23866 40228
rect 23882 40284 23946 40288
rect 23882 40228 23886 40284
rect 23886 40228 23942 40284
rect 23942 40228 23946 40284
rect 23882 40224 23946 40228
rect 23962 40284 24026 40288
rect 23962 40228 23966 40284
rect 23966 40228 24022 40284
rect 24022 40228 24026 40284
rect 23962 40224 24026 40228
rect 27292 40278 27306 40334
rect 27306 40278 27356 40334
rect 27292 40274 27356 40278
rect 31496 40284 31560 40288
rect 31496 40228 31500 40284
rect 31500 40228 31556 40284
rect 31556 40228 31560 40284
rect 31496 40224 31560 40228
rect 31576 40284 31640 40288
rect 31576 40228 31580 40284
rect 31580 40228 31636 40284
rect 31636 40228 31640 40284
rect 31576 40224 31640 40228
rect 31656 40284 31720 40288
rect 31656 40228 31660 40284
rect 31660 40228 31716 40284
rect 31716 40228 31720 40284
rect 31656 40224 31720 40228
rect 31736 40284 31800 40288
rect 31736 40228 31740 40284
rect 31740 40228 31796 40284
rect 31796 40228 31800 40284
rect 31736 40224 31800 40228
rect 14044 40138 14108 40202
rect 28764 40198 28828 40202
rect 28764 40142 28778 40198
rect 28778 40142 28828 40198
rect 28764 40138 28828 40142
rect 8178 40048 8472 40054
rect 8178 39968 8472 40048
rect 12572 40002 12636 40066
rect 16988 40062 17052 40066
rect 16988 40006 17002 40062
rect 17002 40006 17052 40062
rect 16988 40002 17052 40006
rect 8178 39962 8472 39968
rect 2854 39731 2920 39798
rect 30235 39606 30299 39670
rect 28763 39474 28827 39538
rect 31540 39752 31770 39758
rect 31540 39494 31546 39752
rect 31546 39494 31764 39752
rect 31764 39494 31770 39752
rect 31540 39488 31770 39494
rect 27291 39342 27355 39406
rect 25819 39210 25883 39274
rect 24347 39078 24411 39142
rect 22875 38946 22939 39010
rect 21403 38814 21467 38878
rect 18459 38682 18523 38746
rect 16987 38550 17051 38614
rect 15515 38418 15579 38482
rect 14043 38286 14107 38350
rect 12571 38154 12635 38218
rect 11099 38022 11163 38086
rect 9627 37890 9691 37954
rect 7271 37758 7335 37822
rect 5799 37626 5863 37690
rect 4327 37494 4391 37558
rect 5072 31688 5266 31689
rect 5072 31496 5073 31688
rect 5073 31496 5265 31688
rect 5265 31496 5266 31688
rect 5072 31495 5266 31496
rect 26731 31687 26925 31688
rect 26731 31495 26732 31687
rect 26732 31495 26924 31687
rect 26924 31495 26925 31687
rect 26731 31494 26925 31495
rect 5072 29688 5266 29689
rect 5072 29496 5073 29688
rect 5073 29496 5265 29688
rect 5265 29496 5266 29688
rect 5072 29495 5266 29496
rect 26731 29687 26925 29688
rect 26731 29495 26732 29687
rect 26732 29495 26924 29687
rect 26924 29495 26925 29687
rect 26731 29494 26925 29495
rect 5072 27688 5266 27689
rect 5072 27496 5073 27688
rect 5073 27496 5265 27688
rect 5265 27496 5266 27688
rect 5072 27495 5266 27496
rect 26731 27687 26925 27688
rect 26731 27495 26732 27687
rect 26732 27495 26924 27687
rect 26924 27495 26925 27687
rect 26731 27494 26925 27495
rect 5072 25688 5266 25689
rect 5072 25496 5073 25688
rect 5073 25496 5265 25688
rect 5265 25496 5266 25688
rect 5072 25495 5266 25496
rect 26731 25687 26925 25688
rect 26731 25495 26732 25687
rect 26732 25495 26924 25687
rect 26924 25495 26925 25687
rect 26731 25494 26925 25495
rect 5072 23688 5266 23689
rect 5072 23496 5073 23688
rect 5073 23496 5265 23688
rect 5265 23496 5266 23688
rect 5072 23495 5266 23496
rect 26731 23687 26925 23688
rect 26731 23495 26732 23687
rect 26732 23495 26924 23687
rect 26924 23495 26925 23687
rect 26731 23494 26925 23495
rect 5072 21688 5266 21689
rect 5072 21496 5073 21688
rect 5073 21496 5265 21688
rect 5265 21496 5266 21688
rect 5072 21495 5266 21496
rect 26731 21687 26925 21688
rect 26731 21495 26732 21687
rect 26732 21495 26924 21687
rect 26924 21495 26925 21687
rect 26731 21494 26925 21495
rect 5072 19688 5266 19689
rect 5072 19496 5073 19688
rect 5073 19496 5265 19688
rect 5265 19496 5266 19688
rect 5072 19495 5266 19496
rect 26731 19687 26925 19688
rect 26731 19495 26732 19687
rect 26732 19495 26924 19687
rect 26924 19495 26925 19687
rect 26731 19494 26925 19495
rect 5072 17688 5266 17689
rect 5072 17496 5073 17688
rect 5073 17496 5265 17688
rect 5265 17496 5266 17688
rect 5072 17495 5266 17496
rect 26731 17687 26925 17688
rect 26731 17495 26732 17687
rect 26732 17495 26924 17687
rect 26924 17495 26925 17687
rect 26731 17494 26925 17495
rect 5072 15688 5266 15689
rect 5072 15496 5073 15688
rect 5073 15496 5265 15688
rect 5265 15496 5266 15688
rect 5072 15495 5266 15496
rect 26731 15687 26925 15688
rect 26731 15495 26732 15687
rect 26732 15495 26924 15687
rect 26924 15495 26925 15687
rect 26731 15494 26925 15495
rect 5072 13688 5266 13689
rect 5072 13496 5073 13688
rect 5073 13496 5265 13688
rect 5265 13496 5266 13688
rect 5072 13495 5266 13496
rect 26731 13687 26925 13688
rect 26731 13495 26732 13687
rect 26732 13495 26924 13687
rect 26924 13495 26925 13687
rect 26731 13494 26925 13495
rect 5072 11688 5266 11689
rect 5072 11496 5073 11688
rect 5073 11496 5265 11688
rect 5265 11496 5266 11688
rect 5072 11495 5266 11496
rect 26731 11687 26925 11688
rect 26731 11495 26732 11687
rect 26732 11495 26924 11687
rect 26924 11495 26925 11687
rect 26731 11494 26925 11495
rect 5072 9688 5266 9689
rect 5072 9496 5073 9688
rect 5073 9496 5265 9688
rect 5265 9496 5266 9688
rect 5072 9495 5266 9496
rect 26731 9687 26925 9688
rect 26731 9495 26732 9687
rect 26732 9495 26924 9687
rect 26924 9495 26925 9687
rect 26731 9494 26925 9495
rect 5072 7688 5266 7689
rect 5072 7496 5073 7688
rect 5073 7496 5265 7688
rect 5265 7496 5266 7688
rect 5072 7495 5266 7496
rect 26731 7687 26925 7688
rect 26731 7495 26732 7687
rect 26732 7495 26924 7687
rect 26924 7495 26925 7687
rect 26731 7494 26925 7495
rect 5072 5688 5266 5689
rect 5072 5496 5073 5688
rect 5073 5496 5265 5688
rect 5265 5496 5266 5688
rect 5072 5495 5266 5496
rect 26731 5687 26925 5688
rect 26731 5495 26732 5687
rect 26732 5495 26924 5687
rect 26924 5495 26925 5687
rect 26731 5494 26925 5495
rect 5072 3688 5266 3689
rect 5072 3496 5073 3688
rect 5073 3496 5265 3688
rect 5265 3496 5266 3688
rect 5072 3495 5266 3496
rect 26731 3687 26925 3688
rect 26731 3495 26732 3687
rect 26732 3495 26924 3687
rect 26924 3495 26925 3687
rect 26731 3494 26925 3495
rect 5072 1688 5266 1689
rect 5072 1496 5073 1688
rect 5073 1496 5265 1688
rect 5265 1496 5266 1688
rect 5072 1495 5266 1496
rect 26731 1687 26925 1688
rect 26731 1495 26732 1687
rect 26732 1495 26924 1687
rect 26924 1495 26925 1687
rect 26731 1494 26925 1495
<< metal4 >>
rect 798 44555 858 45152
rect 1534 44555 1594 45152
rect 2270 44555 2330 45152
rect 3006 44555 3066 45152
rect 3742 44555 3802 45152
rect 4478 44827 4538 45152
rect 4475 44826 4541 44827
rect 4475 44762 4476 44826
rect 4540 44762 4541 44826
rect 4475 44761 4541 44762
rect 795 44554 861 44555
rect 795 44490 796 44554
rect 860 44490 861 44554
rect 795 44489 861 44490
rect 1531 44554 1597 44555
rect 1531 44490 1532 44554
rect 1596 44490 1597 44554
rect 1531 44489 1597 44490
rect 2267 44554 2333 44555
rect 2267 44490 2268 44554
rect 2332 44490 2333 44554
rect 2267 44489 2333 44490
rect 3003 44554 3069 44555
rect 3003 44490 3004 44554
rect 3068 44490 3069 44554
rect 3003 44489 3069 44490
rect 3739 44554 3805 44555
rect 3739 44490 3740 44554
rect 3804 44490 3805 44554
rect 3739 44489 3805 44490
rect 200 44096 520 44152
rect 200 44032 208 44096
rect 512 44032 520 44096
rect 200 43008 520 44032
rect 200 42944 208 43008
rect 512 42944 520 43008
rect 200 41920 520 42944
rect 200 41856 208 41920
rect 512 41856 520 41920
rect 200 40832 520 41856
rect 4279 44096 4599 44656
rect 5214 44555 5274 45152
rect 5950 44555 6010 45152
rect 5211 44554 5277 44555
rect 5211 44490 5212 44554
rect 5276 44490 5277 44554
rect 5211 44489 5277 44490
rect 5947 44554 6013 44555
rect 5947 44490 5948 44554
rect 6012 44490 6013 44554
rect 5947 44489 6013 44490
rect 4279 44032 4287 44096
rect 4351 44032 4367 44096
rect 4431 44032 4447 44096
rect 4511 44032 4527 44096
rect 4591 44032 4599 44096
rect 4279 43008 4599 44032
rect 4279 42944 4287 43008
rect 4351 42944 4367 43008
rect 4431 42944 4447 43008
rect 4511 42944 4527 43008
rect 4591 42944 4599 43008
rect 4279 41920 4599 42944
rect 4279 41856 4287 41920
rect 4351 41856 4367 41920
rect 4431 41856 4447 41920
rect 4511 41856 4527 41920
rect 4591 41856 4599 41920
rect 1347 41154 1413 41155
rect 1347 41090 1348 41154
rect 1412 41090 1413 41154
rect 1347 41089 1413 41090
rect 2819 41154 2885 41155
rect 2819 41090 2820 41154
rect 2884 41090 2885 41154
rect 2819 41089 2885 41090
rect 200 40768 208 40832
rect 512 40768 520 40832
rect 200 1000 520 40768
rect 1350 40064 1410 41089
rect 2822 40064 2882 41089
rect 4279 40832 4599 41856
rect 6686 41699 6746 45152
rect 7422 42243 7482 45152
rect 8158 44824 8218 45152
rect 7974 44764 8218 44824
rect 7419 42242 7485 42243
rect 7419 42178 7420 42242
rect 7484 42178 7485 42242
rect 7419 42177 7485 42178
rect 7974 42107 8034 44764
rect 8166 44640 8486 44656
rect 8166 44576 8174 44640
rect 8238 44576 8254 44640
rect 8318 44576 8334 44640
rect 8398 44576 8414 44640
rect 8478 44576 8486 44640
rect 8166 43552 8486 44576
rect 8166 43488 8174 43552
rect 8238 43488 8254 43552
rect 8318 43488 8334 43552
rect 8398 43488 8414 43552
rect 8478 43488 8486 43552
rect 8166 42464 8486 43488
rect 8166 42400 8174 42464
rect 8238 42400 8254 42464
rect 8318 42400 8334 42464
rect 8398 42400 8414 42464
rect 8478 42400 8486 42464
rect 7971 42106 8037 42107
rect 7971 42042 7972 42106
rect 8036 42042 8037 42106
rect 7971 42041 8037 42042
rect 6683 41698 6749 41699
rect 6683 41634 6684 41698
rect 6748 41634 6749 41698
rect 6683 41633 6749 41634
rect 4659 41562 4725 41563
rect 4659 41498 4660 41562
rect 4724 41498 4725 41562
rect 4659 41497 4725 41498
rect 4279 40768 4287 40832
rect 4351 40768 4367 40832
rect 4431 40768 4447 40832
rect 4511 40768 4527 40832
rect 4591 40768 4599 40832
rect 4279 40208 4599 40768
rect 4662 40064 4722 41497
rect 8166 41376 8486 42400
rect 8894 41835 8954 45152
rect 9630 44691 9690 45152
rect 9627 44690 9693 44691
rect 9627 44626 9628 44690
rect 9692 44626 9693 44690
rect 9627 44625 9693 44626
rect 10366 41971 10426 45152
rect 10363 41970 10429 41971
rect 10363 41906 10364 41970
rect 10428 41906 10429 41970
rect 10363 41905 10429 41906
rect 8891 41834 8957 41835
rect 8891 41770 8892 41834
rect 8956 41770 8957 41834
rect 8891 41769 8957 41770
rect 11102 41427 11162 45152
rect 8166 41312 8174 41376
rect 8238 41312 8254 41376
rect 8318 41312 8334 41376
rect 8398 41312 8414 41376
rect 8478 41312 8486 41376
rect 11099 41426 11165 41427
rect 11099 41362 11100 41426
rect 11164 41362 11165 41426
rect 11099 41361 11165 41362
rect 5763 41154 5829 41155
rect 5763 41090 5764 41154
rect 5828 41090 5829 41154
rect 5763 41089 5829 41090
rect 7235 41154 7301 41155
rect 7235 41090 7236 41154
rect 7300 41090 7301 41154
rect 7235 41089 7301 41090
rect 1350 40004 1445 40064
rect 2822 40004 2917 40064
rect 1385 39803 1445 40004
rect 2857 39803 2917 40004
rect 4329 40004 4722 40064
rect 5766 40064 5826 41089
rect 7238 40064 7298 41089
rect 8166 40288 8486 41312
rect 11838 41291 11898 45152
rect 12053 44096 12373 44656
rect 12574 44555 12634 45152
rect 12571 44554 12637 44555
rect 12571 44490 12572 44554
rect 12636 44490 12637 44554
rect 12571 44489 12637 44490
rect 12053 44032 12061 44096
rect 12125 44032 12141 44096
rect 12205 44032 12221 44096
rect 12285 44032 12301 44096
rect 12365 44032 12373 44096
rect 12053 43008 12373 44032
rect 12053 42944 12061 43008
rect 12125 42944 12141 43008
rect 12205 42944 12221 43008
rect 12285 42944 12301 43008
rect 12365 42944 12373 43008
rect 12053 41920 12373 42944
rect 13310 42379 13370 45152
rect 14046 43875 14106 45152
rect 14043 43874 14109 43875
rect 14043 43810 14044 43874
rect 14108 43810 14109 43874
rect 14043 43809 14109 43810
rect 14782 43331 14842 45152
rect 15518 44419 15578 45152
rect 16254 44827 16314 45152
rect 16251 44826 16317 44827
rect 16251 44762 16252 44826
rect 16316 44762 16317 44826
rect 16251 44761 16317 44762
rect 15940 44640 16260 44656
rect 15940 44576 15948 44640
rect 16012 44576 16028 44640
rect 16092 44576 16108 44640
rect 16172 44576 16188 44640
rect 16252 44576 16260 44640
rect 15515 44418 15581 44419
rect 15515 44354 15516 44418
rect 15580 44354 15581 44418
rect 15515 44353 15581 44354
rect 15940 43552 16260 44576
rect 16990 44419 17050 45152
rect 17726 44827 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44827 24410 45152
rect 17723 44826 17789 44827
rect 17723 44762 17724 44826
rect 17788 44762 17789 44826
rect 17723 44761 17789 44762
rect 24347 44826 24413 44827
rect 24347 44762 24348 44826
rect 24412 44762 24413 44826
rect 24347 44761 24413 44762
rect 25086 44691 25146 45152
rect 25822 44952 25882 45152
rect 26558 44691 26618 45152
rect 27294 44691 27354 45152
rect 25083 44690 25149 44691
rect 16987 44418 17053 44419
rect 16987 44354 16988 44418
rect 17052 44354 17053 44418
rect 16987 44353 17053 44354
rect 15940 43488 15948 43552
rect 16012 43488 16028 43552
rect 16092 43488 16108 43552
rect 16172 43488 16188 43552
rect 16252 43488 16260 43552
rect 14779 43330 14845 43331
rect 14779 43266 14780 43330
rect 14844 43266 14845 43330
rect 14779 43265 14845 43266
rect 15940 42464 16260 43488
rect 15940 42400 15948 42464
rect 16012 42400 16028 42464
rect 16092 42400 16108 42464
rect 16172 42400 16188 42464
rect 16252 42400 16260 42464
rect 13307 42378 13373 42379
rect 13307 42314 13308 42378
rect 13372 42314 13373 42378
rect 13307 42313 13373 42314
rect 12053 41856 12061 41920
rect 12125 41856 12141 41920
rect 12205 41856 12221 41920
rect 12285 41856 12301 41920
rect 12365 41856 12373 41920
rect 9627 41290 9693 41291
rect 9627 41226 9628 41290
rect 9692 41226 9693 41290
rect 9627 41225 9693 41226
rect 11835 41290 11901 41291
rect 11835 41226 11836 41290
rect 11900 41226 11901 41290
rect 11835 41225 11901 41226
rect 8166 40224 8174 40288
rect 8238 40224 8254 40288
rect 8318 40224 8334 40288
rect 8398 40224 8414 40288
rect 8478 40224 8486 40288
rect 5766 40004 5861 40064
rect 7238 40004 7333 40064
rect 1376 39725 1454 39803
rect 2848 39798 2926 39803
rect 2848 39731 2854 39798
rect 2920 39731 2926 39798
rect 2848 39725 2926 39731
rect 1385 39604 1445 39725
rect 2857 39604 2917 39725
rect 4329 37562 4389 40004
rect 5801 37694 5861 40004
rect 7273 37826 7333 40004
rect 8166 40054 8486 40224
rect 8166 39962 8178 40054
rect 8472 39962 8486 40054
rect 7265 37822 7341 37826
rect 7265 37758 7271 37822
rect 7335 37758 7341 37822
rect 7265 37756 7341 37758
rect 5793 37690 5869 37694
rect 5793 37626 5799 37690
rect 5863 37626 5869 37690
rect 5793 37624 5869 37626
rect 4321 37558 4397 37562
rect 4321 37494 4327 37558
rect 4391 37494 4397 37558
rect 4321 37492 4397 37494
rect 8166 31692 8486 39962
rect 9630 37958 9690 41225
rect 11099 41154 11165 41155
rect 11099 41090 11100 41154
rect 11164 41090 11165 41154
rect 11099 41089 11165 41090
rect 11102 38090 11162 41089
rect 12053 40832 12373 41856
rect 15940 41376 16260 42400
rect 15940 41312 15948 41376
rect 16012 41312 16028 41376
rect 16092 41312 16108 41376
rect 16172 41312 16188 41376
rect 16252 41312 16260 41376
rect 15515 41154 15581 41155
rect 15515 41090 15516 41154
rect 15580 41090 15581 41154
rect 15515 41089 15581 41090
rect 12053 40768 12061 40832
rect 12125 40768 12141 40832
rect 12205 40768 12221 40832
rect 12285 40768 12301 40832
rect 12365 40768 12373 40832
rect 12053 40208 12373 40768
rect 14043 40202 14109 40203
rect 14043 40138 14044 40202
rect 14108 40138 14109 40202
rect 14043 40137 14109 40138
rect 12571 40066 12637 40067
rect 12571 40002 12572 40066
rect 12636 40002 12637 40066
rect 12571 40001 12637 40002
rect 12574 38222 12634 40001
rect 14046 38354 14106 40137
rect 15518 38486 15578 41089
rect 15940 40288 16260 41312
rect 19827 44096 20147 44656
rect 19827 44032 19835 44096
rect 19899 44032 19915 44096
rect 19979 44032 19995 44096
rect 20059 44032 20075 44096
rect 20139 44032 20147 44096
rect 19827 43008 20147 44032
rect 19827 42944 19835 43008
rect 19899 42944 19915 43008
rect 19979 42944 19995 43008
rect 20059 42944 20075 43008
rect 20139 42944 20147 43008
rect 19827 41920 20147 42944
rect 19827 41856 19835 41920
rect 19899 41856 19915 41920
rect 19979 41856 19995 41920
rect 20059 41856 20075 41920
rect 20139 41856 20147 41920
rect 18459 41154 18525 41155
rect 18459 41090 18460 41154
rect 18524 41090 18525 41154
rect 18459 41089 18525 41090
rect 15940 40224 15948 40288
rect 16012 40224 16028 40288
rect 16092 40224 16108 40288
rect 16172 40224 16188 40288
rect 16252 40224 16260 40288
rect 15940 40208 16260 40224
rect 16987 40066 17053 40067
rect 16987 40002 16988 40066
rect 17052 40002 17053 40066
rect 16987 40001 17053 40002
rect 16990 38618 17050 40001
rect 18462 38750 18522 41089
rect 19827 40832 20147 41856
rect 23714 44640 24034 44656
rect 23714 44576 23722 44640
rect 23786 44576 23802 44640
rect 23866 44576 23882 44640
rect 23946 44576 23962 44640
rect 24026 44576 24034 44640
rect 25083 44626 25084 44690
rect 25148 44626 25149 44690
rect 25083 44625 25149 44626
rect 26555 44690 26621 44691
rect 26555 44626 26556 44690
rect 26620 44626 26621 44690
rect 26555 44625 26621 44626
rect 27291 44690 27357 44691
rect 27291 44626 27292 44690
rect 27356 44626 27357 44690
rect 27291 44625 27357 44626
rect 23714 43552 24034 44576
rect 23714 43488 23722 43552
rect 23786 43488 23802 43552
rect 23866 43488 23882 43552
rect 23946 43488 23962 43552
rect 24026 43488 24034 43552
rect 23714 42464 24034 43488
rect 23714 42400 23722 42464
rect 23786 42400 23802 42464
rect 23866 42400 23882 42464
rect 23946 42400 23962 42464
rect 24026 42400 24034 42464
rect 23714 41376 24034 42400
rect 23714 41312 23722 41376
rect 23786 41312 23802 41376
rect 23866 41312 23882 41376
rect 23946 41312 23962 41376
rect 24026 41312 24034 41376
rect 21403 41154 21469 41155
rect 21403 41090 21404 41154
rect 21468 41090 21469 41154
rect 21403 41089 21469 41090
rect 22875 41154 22941 41155
rect 22875 41090 22876 41154
rect 22940 41090 22941 41154
rect 22875 41089 22941 41090
rect 19827 40768 19835 40832
rect 19899 40768 19915 40832
rect 19979 40768 19995 40832
rect 20059 40768 20075 40832
rect 20139 40768 20147 40832
rect 18453 38746 18529 38750
rect 18453 38682 18459 38746
rect 18523 38682 18529 38746
rect 18453 38680 18529 38682
rect 16981 38614 17057 38618
rect 16981 38550 16987 38614
rect 17051 38550 17057 38614
rect 16981 38548 17057 38550
rect 15509 38482 15585 38486
rect 15509 38418 15515 38482
rect 15579 38418 15585 38482
rect 15509 38416 15585 38418
rect 14037 38350 14113 38354
rect 14037 38286 14043 38350
rect 14107 38286 14113 38350
rect 14037 38284 14113 38286
rect 12565 38218 12641 38222
rect 12565 38154 12571 38218
rect 12635 38154 12641 38218
rect 12565 38152 12641 38154
rect 11093 38086 11169 38090
rect 11093 38022 11099 38086
rect 11163 38022 11169 38086
rect 11093 38020 11169 38022
rect 9621 37954 9697 37958
rect 9621 37890 9627 37954
rect 9691 37890 9697 37954
rect 9621 37888 9697 37890
rect 5069 31689 8486 31692
rect 5069 31495 5072 31689
rect 5266 31495 8486 31689
rect 5069 31492 8486 31495
rect 5288 29692 5418 31492
rect 5069 29689 5418 29692
rect 5069 29495 5072 29689
rect 5266 29495 5418 29689
rect 5069 29492 5418 29495
rect 5288 27692 5418 29492
rect 5069 27689 5418 27692
rect 5069 27495 5072 27689
rect 5266 27495 5418 27689
rect 5069 27492 5418 27495
rect 5288 25692 5418 27492
rect 5069 25689 5418 25692
rect 5069 25495 5072 25689
rect 5266 25495 5418 25689
rect 5069 25492 5418 25495
rect 5288 23692 5418 25492
rect 5069 23689 5418 23692
rect 5069 23495 5072 23689
rect 5266 23495 5418 23689
rect 5069 23492 5418 23495
rect 5288 21692 5418 23492
rect 5069 21689 5418 21692
rect 5069 21495 5072 21689
rect 5266 21495 5418 21689
rect 5069 21492 5418 21495
rect 5288 19692 5418 21492
rect 5069 19689 5418 19692
rect 5069 19495 5072 19689
rect 5266 19495 5418 19689
rect 5069 19492 5418 19495
rect 5288 17692 5418 19492
rect 5069 17689 5418 17692
rect 5069 17495 5072 17689
rect 5266 17495 5418 17689
rect 5069 17492 5418 17495
rect 5288 15692 5418 17492
rect 5069 15689 5418 15692
rect 5069 15495 5072 15689
rect 5266 15495 5418 15689
rect 5069 15492 5418 15495
rect 5288 13692 5418 15492
rect 5069 13689 5418 13692
rect 5069 13495 5072 13689
rect 5266 13495 5418 13689
rect 5069 13492 5418 13495
rect 5288 11692 5418 13492
rect 5069 11689 5418 11692
rect 5069 11495 5072 11689
rect 5266 11495 5418 11689
rect 5069 11492 5418 11495
rect 5288 9692 5418 11492
rect 5069 9689 5418 9692
rect 5069 9495 5072 9689
rect 5266 9495 5418 9689
rect 5069 9492 5418 9495
rect 5288 7692 5418 9492
rect 5069 7689 5418 7692
rect 5069 7495 5072 7689
rect 5266 7495 5418 7689
rect 5069 7492 5418 7495
rect 5288 5692 5418 7492
rect 5069 5689 5418 5692
rect 5069 5495 5072 5689
rect 5266 5495 5418 5689
rect 5069 5492 5418 5495
rect 5288 3692 5418 5492
rect 5069 3689 5418 3692
rect 5069 3495 5072 3689
rect 5266 3495 5418 3689
rect 5069 3492 5418 3495
rect 5288 1692 5418 3492
rect 8166 1692 8486 31492
rect 5069 1689 8486 1692
rect 5069 1495 5072 1689
rect 5266 1495 8486 1689
rect 5069 1492 8486 1495
rect 5288 1491 5418 1492
rect 8166 1000 8486 1492
rect 19827 31691 20147 40768
rect 21406 38882 21466 41089
rect 22878 39014 22938 41089
rect 23714 40288 24034 41312
rect 27601 44096 27921 44656
rect 28030 44147 28090 45152
rect 27601 44032 27609 44096
rect 27673 44032 27689 44096
rect 27753 44032 27769 44096
rect 27833 44032 27849 44096
rect 27913 44032 27921 44096
rect 28027 44146 28093 44147
rect 28027 44082 28028 44146
rect 28092 44082 28093 44146
rect 28027 44081 28093 44082
rect 27601 43008 27921 44032
rect 28766 43875 28826 45152
rect 29502 44147 29562 45152
rect 29499 44146 29565 44147
rect 29499 44082 29500 44146
rect 29564 44082 29565 44146
rect 29499 44081 29565 44082
rect 28763 43874 28829 43875
rect 28763 43810 28764 43874
rect 28828 43810 28829 43874
rect 28763 43809 28829 43810
rect 27601 42944 27609 43008
rect 27673 42944 27689 43008
rect 27753 42944 27769 43008
rect 27833 42944 27849 43008
rect 27913 42944 27921 43008
rect 27601 41920 27921 42944
rect 30238 42243 30298 45152
rect 30974 44011 31034 45152
rect 31710 44824 31770 45152
rect 31342 44764 31770 44824
rect 30971 44010 31037 44011
rect 30971 43946 30972 44010
rect 31036 43946 31037 44010
rect 30971 43945 31037 43946
rect 30235 42242 30301 42243
rect 30235 42178 30236 42242
rect 30300 42178 30301 42242
rect 30235 42177 30301 42178
rect 27601 41856 27609 41920
rect 27673 41856 27689 41920
rect 27753 41856 27769 41920
rect 27833 41856 27849 41920
rect 27913 41856 27921 41920
rect 24347 41154 24413 41155
rect 24347 41090 24348 41154
rect 24412 41090 24413 41154
rect 24347 41089 24413 41090
rect 25819 41154 25885 41155
rect 25819 41090 25820 41154
rect 25884 41090 25885 41154
rect 25819 41089 25885 41090
rect 23714 40224 23722 40288
rect 23786 40224 23802 40288
rect 23866 40224 23882 40288
rect 23946 40224 23962 40288
rect 24026 40224 24034 40288
rect 23714 40208 24034 40224
rect 24350 39146 24410 41089
rect 25822 39278 25882 41089
rect 27601 40832 27921 41856
rect 31342 41835 31402 44764
rect 31488 44640 31808 44656
rect 31488 44576 31496 44640
rect 31560 44576 31576 44640
rect 31640 44576 31656 44640
rect 31720 44576 31736 44640
rect 31800 44576 31808 44640
rect 31488 43552 31808 44576
rect 31488 43488 31496 43552
rect 31560 43488 31576 43552
rect 31640 43488 31656 43552
rect 31720 43488 31736 43552
rect 31800 43488 31808 43552
rect 31488 42464 31808 43488
rect 31488 42400 31496 42464
rect 31560 42400 31576 42464
rect 31640 42400 31656 42464
rect 31720 42400 31736 42464
rect 31800 42400 31808 42464
rect 31339 41834 31405 41835
rect 31339 41770 31340 41834
rect 31404 41770 31405 41834
rect 31339 41769 31405 41770
rect 31488 41376 31808 42400
rect 31488 41312 31496 41376
rect 31560 41312 31576 41376
rect 31640 41312 31656 41376
rect 31720 41312 31736 41376
rect 31800 41312 31808 41376
rect 30235 41154 30301 41155
rect 30235 41090 30236 41154
rect 30300 41090 30301 41154
rect 30235 41089 30301 41090
rect 27601 40768 27609 40832
rect 27673 40768 27689 40832
rect 27753 40768 27769 40832
rect 27833 40768 27849 40832
rect 27913 40768 27921 40832
rect 27291 40338 27357 40339
rect 27291 40274 27292 40338
rect 27356 40274 27357 40338
rect 27291 40273 27357 40274
rect 27294 39410 27354 40273
rect 27601 40208 27921 40768
rect 28763 40202 28829 40203
rect 28763 40138 28764 40202
rect 28828 40138 28829 40202
rect 28763 40137 28829 40138
rect 28766 39542 28826 40137
rect 30238 39674 30298 41089
rect 31488 40288 31808 41312
rect 31488 40224 31496 40288
rect 31560 40224 31576 40288
rect 31640 40224 31656 40288
rect 31720 40224 31736 40288
rect 31800 40224 31808 40288
rect 31488 39758 31808 40224
rect 30229 39670 30305 39674
rect 30229 39606 30235 39670
rect 30299 39606 30305 39670
rect 30229 39604 30305 39606
rect 28757 39538 28833 39542
rect 28757 39474 28763 39538
rect 28827 39474 28833 39538
rect 28757 39472 28833 39474
rect 31488 39488 31540 39758
rect 31770 39488 31808 39758
rect 27285 39406 27361 39410
rect 27285 39342 27291 39406
rect 27355 39342 27361 39406
rect 27285 39340 27361 39342
rect 25813 39274 25889 39278
rect 25813 39210 25819 39274
rect 25883 39210 25889 39274
rect 25813 39208 25889 39210
rect 24341 39142 24417 39146
rect 24341 39078 24347 39142
rect 24411 39078 24417 39142
rect 24341 39076 24417 39078
rect 22869 39010 22945 39014
rect 22869 38946 22875 39010
rect 22939 38946 22945 39010
rect 22869 38944 22945 38946
rect 21397 38878 21473 38882
rect 21397 38814 21403 38878
rect 21467 38814 21473 38878
rect 21397 38812 21473 38814
rect 19827 31688 26928 31691
rect 19827 31494 26731 31688
rect 26925 31494 26928 31688
rect 19827 31491 26928 31494
rect 19827 1691 20147 31491
rect 26578 29691 26708 31491
rect 26578 29688 26928 29691
rect 26578 29494 26731 29688
rect 26925 29494 26928 29688
rect 26578 29491 26928 29494
rect 26578 27691 26708 29491
rect 26578 27688 26928 27691
rect 26578 27494 26731 27688
rect 26925 27494 26928 27688
rect 26578 27491 26928 27494
rect 26578 25691 26708 27491
rect 26578 25688 26928 25691
rect 26578 25494 26731 25688
rect 26925 25494 26928 25688
rect 26578 25491 26928 25494
rect 26578 23691 26708 25491
rect 26578 23688 26928 23691
rect 26578 23494 26731 23688
rect 26925 23494 26928 23688
rect 26578 23491 26928 23494
rect 26578 21691 26708 23491
rect 26578 21688 26928 21691
rect 26578 21494 26731 21688
rect 26925 21494 26928 21688
rect 26578 21491 26928 21494
rect 26578 19691 26708 21491
rect 26578 19688 26928 19691
rect 26578 19494 26731 19688
rect 26925 19494 26928 19688
rect 26578 19491 26928 19494
rect 26578 17691 26708 19491
rect 26578 17688 26928 17691
rect 26578 17494 26731 17688
rect 26925 17494 26928 17688
rect 26578 17491 26928 17494
rect 26578 15691 26708 17491
rect 26578 15688 26928 15691
rect 26578 15494 26731 15688
rect 26925 15494 26928 15688
rect 26578 15491 26928 15494
rect 26578 13691 26708 15491
rect 26578 13688 26928 13691
rect 26578 13494 26731 13688
rect 26925 13494 26928 13688
rect 26578 13491 26928 13494
rect 26578 11691 26708 13491
rect 26578 11688 26928 11691
rect 26578 11494 26731 11688
rect 26925 11494 26928 11688
rect 26578 11491 26928 11494
rect 26578 9691 26708 11491
rect 26578 9688 26928 9691
rect 26578 9494 26731 9688
rect 26925 9494 26928 9688
rect 26578 9491 26928 9494
rect 26578 7691 26708 9491
rect 26578 7688 26928 7691
rect 26578 7494 26731 7688
rect 26925 7494 26928 7688
rect 26578 7491 26928 7494
rect 26578 5691 26708 7491
rect 26578 5688 26928 5691
rect 26578 5494 26731 5688
rect 26925 5494 26928 5688
rect 26578 5491 26928 5494
rect 26578 3691 26708 5491
rect 26578 3688 26928 3691
rect 26578 3494 26731 3688
rect 26925 3494 26928 3688
rect 26578 3491 26928 3494
rect 26578 1691 26708 3491
rect 19827 1688 26928 1691
rect 19827 1494 26731 1688
rect 26925 1494 26928 1688
rect 19827 1491 26928 1494
rect 19827 1000 20147 1491
rect 31488 1000 31808 39488
rect 370 0 550 200
rect 4786 0 4966 200
rect 9202 0 9382 200
rect 13618 0 13798 200
rect 18034 0 18214 200
rect 22450 0 22630 200
rect 26866 0 27046 200
rect 31282 0 31462 200
use sky130_fd_sc_hd__clkbuf_8  _059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 13156 0 -1 43520
box -38 -48 1050 592
use sky130_fd_sc_hd__or2b_1  _060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 25392 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 26956 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 25300 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 23000 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 15272 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _065_
timestamp 1707688321
transform -1 0 18584 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _066_
timestamp 1707688321
transform 1 0 22724 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _067_
timestamp 1707688321
transform -1 0 16008 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _068_
timestamp 1707688321
transform 1 0 22724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _069_
timestamp 1707688321
transform 1 0 18676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _070_
timestamp 1707688321
transform 1 0 22724 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _071_
timestamp 1707688321
transform 1 0 19412 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 22632 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 17388 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 16928 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 16928 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _076_
timestamp 1707688321
transform 1 0 16928 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _077_
timestamp 1707688321
transform 1 0 14720 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _078_
timestamp 1707688321
transform 1 0 15180 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 13984 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 14352 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _081_
timestamp 1707688321
transform -1 0 12420 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_4  _082_
timestamp 1707688321
transform 1 0 12972 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _083_
timestamp 1707688321
transform -1 0 13340 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 12972 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 11684 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_1  _086_
timestamp 1707688321
transform -1 0 12880 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _087_
timestamp 1707688321
transform -1 0 11408 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 14904 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 11408 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _090_
timestamp 1707688321
transform 1 0 12880 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _091_
timestamp 1707688321
transform 1 0 16284 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _092_
timestamp 1707688321
transform -1 0 18216 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _093_
timestamp 1707688321
transform -1 0 16376 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _094_
timestamp 1707688321
transform -1 0 14904 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _095_
timestamp 1707688321
transform -1 0 14352 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 14904 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _097_
timestamp 1707688321
transform -1 0 14076 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _098_
timestamp 1707688321
transform -1 0 13248 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _099_
timestamp 1707688321
transform -1 0 11960 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1707688321
transform -1 0 13800 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 15364 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__nor3_4  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 13708 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1707688321
transform 1 0 20148 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 13156 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 6808 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _106_
timestamp 1707688321
transform -1 0 16560 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1707688321
transform -1 0 8280 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _108_
timestamp 1707688321
transform -1 0 12512 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _109_
timestamp 1707688321
transform 1 0 11684 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _110_
timestamp 1707688321
transform -1 0 15824 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _111_
timestamp 1707688321
transform -1 0 15180 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _112_
timestamp 1707688321
transform -1 0 16008 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _113_
timestamp 1707688321
transform 1 0 15364 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1707688321
transform 1 0 16100 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _115_
timestamp 1707688321
transform 1 0 16928 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1707688321
transform 1 0 17756 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _117_
timestamp 1707688321
transform 1 0 19228 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1707688321
transform 1 0 20240 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _119_
timestamp 1707688321
transform 1 0 20516 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1707688321
transform 1 0 21988 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 14076 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1707688321
transform 1 0 23460 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _123_
timestamp 1707688321
transform 1 0 19412 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _124_
timestamp 1707688321
transform 1 0 20608 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _125_
timestamp 1707688321
transform -1 0 22264 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _126_
timestamp 1707688321
transform -1 0 21988 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _127_
timestamp 1707688321
transform 1 0 17940 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _128_
timestamp 1707688321
transform 1 0 19136 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 24380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 23460 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1707688321
transform 1 0 21988 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _132_
timestamp 1707688321
transform 1 0 21252 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _133_
timestamp 1707688321
transform 1 0 24564 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1707688321
transform 1 0 26404 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _135_
timestamp 1707688321
transform 1 0 25392 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 30636 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1707688321
transform 1 0 30452 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1707688321
transform -1 0 29808 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1707688321
transform 1 0 29256 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1707688321
transform -1 0 28888 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1707688321
transform 1 0 29164 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1707688321
transform 1 0 26864 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1707688321
transform 1 0 26864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144__1
timestamp 1707688321
transform -1 0 24104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1707688321
transform 1 0 20424 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1707688321
transform 1 0 19872 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147__2
timestamp 1707688321
transform 1 0 19228 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__3
timestamp 1707688321
transform 1 0 14996 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149__4
timestamp 1707688321
transform 1 0 15732 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150__5
timestamp 1707688321
transform 1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 23000 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _152_
timestamp 1707688321
transform 1 0 24380 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 19320 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _154_
timestamp 1707688321
transform 1 0 29440 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _155_
timestamp 1707688321
transform 1 0 28980 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _156_
timestamp 1707688321
transform -1 0 28888 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _157_
timestamp 1707688321
transform 1 0 26588 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _158_
timestamp 1707688321
transform 1 0 24472 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _159_
timestamp 1707688321
transform 1 0 24288 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _160_
timestamp 1707688321
transform 1 0 23552 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 19688 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_2  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 19136 0 -1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _163_
timestamp 1707688321
transform 1 0 15824 0 1 43520
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _164_
timestamp 1707688321
transform 1 0 16100 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _165_
timestamp 1707688321
transform 1 0 11684 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _166_
timestamp 1707688321
transform 1 0 20056 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _176_
timestamp 1707688321
transform -1 0 4600 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _177_
timestamp 1707688321
transform -1 0 2392 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _178_
timestamp 1707688321
transform -1 0 14352 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  amux_ctrl.async_and3.genblk1.genblk1.genblk1.and3_2_dont_touch $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 22356 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  amux_ctrl.async_nor2.genblk1.genblk1.genblk1.nor2_2_dont_touch $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 22724 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  amux_ctrl.por_0_dfxtp_2.genblk1.genblk1.genblk1.dfxtp_2_dont_touch
timestamp 1707688321
transform 1 0 3864 0 1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dlygate4sd3_1  amux_ctrl.por_0_dlygate4sd3_1.genblk1.genblk1.dlygate4sd3_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5980 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  amux_ctrl.por_1_dfxtp_2.genblk1.genblk1.genblk1.dfxtp_2_dont_touch
timestamp 1707688321
transform -1 0 3956 0 -1 41344
box -38 -48 1602 592
use sky130_fd_sc_hd__dlygate4sd3_1  amux_ctrl.por_1_dlygate4sd3_1.genblk1.genblk1.dlygate4sd3_1
timestamp 1707688321
transform 1 0 3404 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  amux_ctrl.por_2_dfxtp_1.genblk1.genblk1.dfxtp_1_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 2392 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  amux_ctrl.por_2_dfxtp_1.genblk1.genblk1.dfxtp_1
timestamp 1707688321
transform -1 0 3312 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  amux_ctrl.por_2_dlygate4sd3_1.genblk1.genblk1.dlygate4sd3_1
timestamp 1707688321
transform 1 0 2392 0 1 41344
box -38 -48 774 592
use tt07_1v8_analog_io_2wire  tt07_1v8_analog_io_2wire_0_0
timestamp 1717291860
transform 1 0 0 0 1 0
box 1770 0 31472 1200
use sky130_fd_sc_hd__buf_4  buf_oa_ena.genblk1.genblk1.genblk1.genblk1.buf_4_dont_touch $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 30544 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform -1 0 18216 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1707688321
transform -1 0 13156 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1707688321
transform 1 0 21436 0 -1 43520
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 828 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1707688321
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3036 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1707688321
transform 1 0 3220 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1707688321
transform 1 0 4324 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 5428 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1707688321
transform 1 0 5796 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1707688321
transform 1 0 6900 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1707688321
transform 1 0 8004 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1707688321
transform 1 0 8372 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1707688321
transform 1 0 9476 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1707688321
transform 1 0 10580 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1707688321
transform 1 0 10948 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 12052 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_131
timestamp 1707688321
transform 1 0 12604 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1707688321
transform 1 0 13156 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1707688321
transform 1 0 13524 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 14628 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1717249547
transform 1 0 15824 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_173
timestamp 1707688321
transform 1 0 16468 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_185 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 17572 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1707688321
transform 1 0 18308 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1707688321
transform 1 0 18676 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1707688321
transform 1 0 19780 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1707688321
transform 1 0 20884 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1707688321
transform 1 0 21252 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1707688321
transform 1 0 22356 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1707688321
transform 1 0 23460 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1707688321
transform 1 0 23828 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1707688321
transform 1 0 24932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1707688321
transform 1 0 26036 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1707688321
transform 1 0 26404 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1707688321
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1707688321
transform 1 0 28612 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1707688321
transform 1 0 28980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1707688321
transform 1 0 30084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_333
timestamp 1717249547
transform 1 0 31188 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1707688321
transform 1 0 828 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_15
timestamp 1707688321
transform 1 0 1932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_37
timestamp 1707688321
transform 1 0 3956 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_44
timestamp 1707688321
transform 1 0 4600 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1707688321
transform 1 0 5796 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1707688321
transform 1 0 6348 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_68
timestamp 1707688321
transform 1 0 6808 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_84
timestamp 1707688321
transform 1 0 8280 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_96
timestamp 1707688321
transform 1 0 9384 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_108
timestamp 1707688321
transform 1 0 10488 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1707688321
transform 1 0 10948 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_191
timestamp 1707688321
transform 1 0 18124 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_199
timestamp 1707688321
transform 1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_208
timestamp 1707688321
transform 1 0 19688 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 1717249547
transform 1 0 21252 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1707688321
transform 1 0 22356 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_252
timestamp 1707688321
transform 1 0 23736 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_264
timestamp 1707688321
transform 1 0 24840 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_276
timestamp 1707688321
transform 1 0 25944 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1707688321
transform 1 0 26404 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1707688321
transform 1 0 27508 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1707688321
transform 1 0 28612 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_317
timestamp 1707688321
transform 1 0 29716 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_326
timestamp 1707688321
transform 1 0 30544 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_334
timestamp 1707688321
transform 1 0 31280 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1707688321
transform 1 0 828 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_15
timestamp 1717249547
transform 1 0 1932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 1707688321
transform 1 0 3220 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 1707688321
transform 1 0 3772 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_53
timestamp 1707688321
transform 1 0 5428 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_67
timestamp 1707688321
transform 1 0 6716 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_79
timestamp 1707688321
transform 1 0 7820 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1707688321
transform 1 0 8188 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1707688321
transform 1 0 8372 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1707688321
transform 1 0 9476 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1707688321
transform 1 0 10580 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1707688321
transform 1 0 13340 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_144
timestamp 1707688321
transform 1 0 13800 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_166
timestamp 1707688321
transform 1 0 15824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_183
timestamp 1707688321
transform 1 0 17388 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1717249547
transform 1 0 18400 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_197
timestamp 1707688321
transform 1 0 18676 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1707688321
transform 1 0 22724 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1707688321
transform 1 0 23460 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1707688321
transform 1 0 23828 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_265
timestamp 1707688321
transform 1 0 24932 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_269
timestamp 1707688321
transform 1 0 25300 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_276
timestamp 1707688321
transform 1 0 25944 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_288
timestamp 1707688321
transform 1 0 27048 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_300
timestamp 1707688321
transform 1 0 28152 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1707688321
transform 1 0 28980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1707688321
transform 1 0 30084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_333
timestamp 1717249547
transform 1 0 31188 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3
timestamp 1707688321
transform 1 0 828 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_11
timestamp 1707688321
transform 1 0 1564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_30
timestamp 1707688321
transform 1 0 3312 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1707688321
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1707688321
transform 1 0 5244 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1707688321
transform 1 0 5612 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1707688321
transform 1 0 5796 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1707688321
transform 1 0 6900 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1707688321
transform 1 0 8004 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1707688321
transform 1 0 9108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1707688321
transform 1 0 10212 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1707688321
transform 1 0 10764 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 1707688321
transform 1 0 10948 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_117
timestamp 1707688321
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_144
timestamp 1707688321
transform 1 0 13800 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_155
timestamp 1707688321
transform 1 0 14812 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_183
timestamp 1707688321
transform 1 0 17388 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_195
timestamp 1707688321
transform 1 0 18492 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_203
timestamp 1717249547
transform 1 0 19228 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_240
timestamp 1707688321
transform 1 0 22632 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_249
timestamp 1707688321
transform 1 0 23460 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_257
timestamp 1707688321
transform 1 0 24196 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_276
timestamp 1707688321
transform 1 0 25944 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_289
timestamp 1707688321
transform 1 0 27140 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_301
timestamp 1707688321
transform 1 0 28244 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_313
timestamp 1707688321
transform 1 0 29348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_325
timestamp 1707688321
transform 1 0 30452 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_333
timestamp 1717249547
transform 1 0 31188 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1707688321
transform 1 0 828 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1707688321
transform 1 0 1932 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1707688321
transform 1 0 3036 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1707688321
transform 1 0 3220 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1707688321
transform 1 0 4324 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1707688321
transform 1 0 5428 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1707688321
transform 1 0 6532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1707688321
transform 1 0 7636 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1707688321
transform 1 0 8188 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1707688321
transform 1 0 8372 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1707688321
transform 1 0 9476 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_109
timestamp 1707688321
transform 1 0 10580 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_150
timestamp 1707688321
transform 1 0 14352 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1707688321
transform 1 0 18676 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_209
timestamp 1707688321
transform 1 0 19780 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_215
timestamp 1707688321
transform 1 0 20332 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_287
timestamp 1707688321
transform 1 0 26956 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_295
timestamp 1707688321
transform 1 0 27692 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1717249547
transform 1 0 28704 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_315
timestamp 1707688321
transform 1 0 29532 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_323
timestamp 1717249547
transform 1 0 30268 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_328
timestamp 1707688321
transform 1 0 30728 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_334
timestamp 1707688321
transform 1 0 31280 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1707688321
transform 1 0 828 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1707688321
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1707688321
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1707688321
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1707688321
transform 1 0 5244 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1707688321
transform 1 0 5612 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1707688321
transform 1 0 5796 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1707688321
transform 1 0 6900 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1707688321
transform 1 0 8004 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1707688321
transform 1 0 9108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1707688321
transform 1 0 10212 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1707688321
transform 1 0 10764 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_113
timestamp 1707688321
transform 1 0 10948 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_163
timestamp 1717249547
transform 1 0 15548 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_202
timestamp 1717249547
transform 1 0 19136 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_225
timestamp 1717249547
transform 1 0 21252 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_247
timestamp 1707688321
transform 1 0 23276 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_269
timestamp 1707688321
transform 1 0 25300 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_284
timestamp 1717249547
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_289
timestamp 1707688321
transform 1 0 27140 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_333
timestamp 1717249547
transform 1 0 31188 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1707688321
transform 1 0 828 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1707688321
transform 1 0 1932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1707688321
transform 1 0 3036 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1707688321
transform 1 0 3220 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1707688321
transform 1 0 4324 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1707688321
transform 1 0 5428 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1707688321
transform 1 0 6532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1707688321
transform 1 0 7636 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1707688321
transform 1 0 8188 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1707688321
transform 1 0 8372 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1707688321
transform 1 0 9476 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_109
timestamp 1707688321
transform 1 0 10580 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1707688321
transform 1 0 13156 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_156
timestamp 1707688321
transform 1 0 14904 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_192
timestamp 1707688321
transform 1 0 18216 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_211
timestamp 1707688321
transform 1 0 19964 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_256
timestamp 1717249547
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_274
timestamp 1707688321
transform 1 0 25760 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_282
timestamp 1707688321
transform 1 0 26496 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_325
timestamp 1707688321
transform 1 0 30452 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_334
timestamp 1707688321
transform 1 0 31280 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_6
timestamp 1707688321
transform 1 0 1104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_10
timestamp 1707688321
transform 1 0 1472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_14
timestamp 1707688321
transform 1 0 1840 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_18
timestamp 1707688321
transform 1 0 2208 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_22
timestamp 1707688321
transform 1 0 2576 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_32
timestamp 1707688321
transform 1 0 3496 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_38
timestamp 1707688321
transform 1 0 4048 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_42
timestamp 1707688321
transform 1 0 4416 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_46
timestamp 1707688321
transform 1 0 4784 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_50
timestamp 1707688321
transform 1 0 5152 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1717249547
transform 1 0 5520 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1717249547
transform 1 0 5796 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_62
timestamp 1707688321
transform 1 0 6256 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_74
timestamp 1707688321
transform 1 0 7360 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_82
timestamp 1717249547
transform 1 0 8096 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_85
timestamp 1707688321
transform 1 0 8372 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_97
timestamp 1707688321
transform 1 0 9476 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_109
timestamp 1707688321
transform 1 0 10580 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1707688321
transform 1 0 10948 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1707688321
transform 1 0 11500 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_129
timestamp 1707688321
transform 1 0 12420 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_138
timestamp 1717249547
transform 1 0 13248 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_150
timestamp 1707688321
transform 1 0 14352 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1717249547
transform 1 0 16100 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_180
timestamp 1707688321
transform 1 0 17112 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_191
timestamp 1707688321
transform 1 0 18124 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_195
timestamp 1707688321
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_206
timestamp 1707688321
transform 1 0 19504 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_218
timestamp 1707688321
transform 1 0 20608 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_236
timestamp 1707688321
transform 1 0 22264 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_240
timestamp 1707688321
transform 1 0 22632 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp 1707688321
transform 1 0 23460 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_253
timestamp 1707688321
transform 1 0 23828 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_272
timestamp 1707688321
transform 1 0 25576 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1717249547
transform 1 0 26404 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_306
timestamp 1717249547
transform 1 0 28704 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1707688321
transform -1 0 26588 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1707688321
transform -1 0 21988 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1707688321
transform -1 0 22724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1707688321
transform -1 0 21988 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1707688321
transform -1 0 27140 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1707688321
transform 1 0 18676 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1707688321
transform 1 0 17388 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1707688321
transform -1 0 28428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1707688321
transform 1 0 27968 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1707688321
transform -1 0 31372 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1707688321
transform -1 0 31280 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1707688321
transform 1 0 30912 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1707688321
transform -1 0 29256 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1707688321
transform 1 0 28888 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1707688321
transform 1 0 28428 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1707688321
transform 1 0 26588 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1707688321
transform 1 0 25300 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1707688321
transform 1 0 25024 0 -1 44608
box -38 -48 314 592
use my_transmission_gate_in_00  my_transmission_gate_in_00 my_transmission_gate_in/00
timestamp 1717265471
transform 1 0 200 0 1 1200
box 0 0 5070 2100
use my_transmission_gate_in_01  my_transmission_gate_in_01 my_transmission_gate_in/01
timestamp 1717265471
transform 1 0 200 0 1 3200
box 0 0 5070 2100
use my_transmission_gate_in_02  my_transmission_gate_in_02 my_transmission_gate_in/02
timestamp 1717265471
transform 1 0 200 0 1 5200
box 0 0 5070 2100
use my_transmission_gate_in_03  my_transmission_gate_in_03 my_transmission_gate_in/03
timestamp 1717265471
transform 1 0 200 0 1 7200
box 0 0 5070 2100
use my_transmission_gate_in_04  my_transmission_gate_in_04 my_transmission_gate_in/04
timestamp 1717265471
transform 1 0 200 0 1 9200
box 0 0 5070 2100
use my_transmission_gate_in_05  my_transmission_gate_in_05 my_transmission_gate_in/05
timestamp 1717265471
transform 1 0 200 0 1 11200
box 0 0 5070 2100
use my_transmission_gate_in_06  my_transmission_gate_in_06 my_transmission_gate_in/06
timestamp 1717265471
transform 1 0 200 0 1 13200
box 0 0 5070 2100
use my_transmission_gate_in_07  my_transmission_gate_in_07 my_transmission_gate_in/07
timestamp 1717265471
transform 1 0 200 0 1 15200
box 0 0 5070 2100
use my_transmission_gate_in_08  my_transmission_gate_in_08 my_transmission_gate_in/08
timestamp 1717265471
transform 1 0 200 0 1 17200
box 0 0 5070 2100
use my_transmission_gate_in_09  my_transmission_gate_in_09 my_transmission_gate_in/09
timestamp 1717265471
transform 1 0 200 0 1 19200
box 0 0 5070 2100
use my_transmission_gate_in_10  my_transmission_gate_in_10 my_transmission_gate_in/10
timestamp 1717265471
transform 1 0 200 0 1 21200
box 0 0 5070 2100
use my_transmission_gate_in_11  my_transmission_gate_in_11 my_transmission_gate_in/11
timestamp 1717265471
transform 1 0 200 0 1 23200
box 0 0 5070 2100
use my_transmission_gate_in_12  my_transmission_gate_in_12 my_transmission_gate_in/12
timestamp 1717265471
transform 1 0 200 0 1 25200
box 0 0 5070 2100
use my_transmission_gate_in_13  my_transmission_gate_in_13 my_transmission_gate_in/13
timestamp 1717265471
transform 1 0 200 0 1 27200
box 0 0 5070 2100
use my_transmission_gate_in_14  my_transmission_gate_in_14 my_transmission_gate_in/14
timestamp 1717265471
transform 1 0 200 0 1 29200
box 0 0 5070 2100
use my_transmission_gate_in_15  my_transmission_gate_in_15 my_transmission_gate_in/15
timestamp 1717265471
transform 1 0 200 0 1 31200
box 0 0 5070 2100
use my_transmission_gate_out_00  my_transmission_gate_out_00 my_transmission_gate_out/00
timestamp 1717289656
transform 1 0 26728 0 1 1198
box 0 0 5080 2100
use my_transmission_gate_out_01  my_transmission_gate_out_01 my_transmission_gate_out/01
timestamp 1717261669
transform 1 0 26728 0 1 3198
box 0 0 5080 2100
use my_transmission_gate_out_02  my_transmission_gate_out_02 my_transmission_gate_out/02
timestamp 1717261669
transform 1 0 26728 0 1 5198
box 0 0 5080 2100
use my_transmission_gate_out_03  my_transmission_gate_out_03 my_transmission_gate_out/03
timestamp 1717261669
transform 1 0 26728 0 1 7198
box 0 0 5080 2100
use my_transmission_gate_out_04  my_transmission_gate_out_04 my_transmission_gate_out/04
timestamp 1717261669
transform 1 0 26728 0 1 9198
box 0 0 5080 2100
use my_transmission_gate_out_05  my_transmission_gate_out_05 my_transmission_gate_out/05
timestamp 1717261669
transform 1 0 26728 0 1 11198
box 0 0 5080 2100
use my_transmission_gate_out_06  my_transmission_gate_out_06 my_transmission_gate_out/06
timestamp 1717261669
transform 1 0 26728 0 1 13198
box 0 0 5080 2100
use my_transmission_gate_out_07  my_transmission_gate_out_07 my_transmission_gate_out/07
timestamp 1717261669
transform 1 0 26728 0 1 15198
box 0 0 5080 2100
use my_transmission_gate_out_08  my_transmission_gate_out_08 my_transmission_gate_out/08
timestamp 1717261669
transform 1 0 26728 0 1 17198
box 0 0 5080 2100
use my_transmission_gate_out_09  my_transmission_gate_out_09 my_transmission_gate_out/09
timestamp 1717261669
transform 1 0 26728 0 1 19198
box 0 0 5080 2100
use my_transmission_gate_out_10  my_transmission_gate_out_10 my_transmission_gate_out/10
timestamp 1717260747
transform 1 0 26728 0 1 21198
box 0 0 5080 2100
use my_transmission_gate_out_11  my_transmission_gate_out_11 my_transmission_gate_out/11
timestamp 1717260747
transform 1 0 26728 0 1 23198
box 0 0 5080 2100
use my_transmission_gate_out_12  my_transmission_gate_out_12 my_transmission_gate_out/12
timestamp 1717260747
transform 1 0 26728 0 1 25198
box 0 0 5080 2100
use my_transmission_gate_out_13  my_transmission_gate_out_13 my_transmission_gate_out/13
timestamp 1717260747
transform 1 0 26728 0 1 27198
box 0 0 5080 2100
use my_transmission_gate_out_14  my_transmission_gate_out_14 my_transmission_gate_out/14
timestamp 1717260013
transform 1 0 26728 0 1 29198
box 0 0 5080 2100
use my_transmission_gate_out_15  my_transmission_gate_out_15 my_transmission_gate_out/15
timestamp 1717260013
transform 1 0 26728 0 1 31198
box 0 0 5080 2100
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_8
timestamp 1707688321
transform 1 0 552 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1707688321
transform -1 0 31648 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_9
timestamp 1707688321
transform 1 0 552 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1707688321
transform -1 0 31648 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_10
timestamp 1707688321
transform 1 0 552 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1707688321
transform -1 0 31648 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_11
timestamp 1707688321
transform 1 0 552 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1707688321
transform -1 0 31648 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_12
timestamp 1707688321
transform 1 0 552 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1707688321
transform -1 0 31648 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_13
timestamp 1707688321
transform 1 0 552 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1707688321
transform -1 0 31648 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_14
timestamp 1707688321
transform 1 0 552 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1707688321
transform -1 0 31648 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_15
timestamp 1707688321
transform 1 0 552 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1707688321
transform -1 0 31648 0 -1 44608
box -38 -48 314 592
use sky130_fd_pr__res_xhigh_po_0p35_PYW3KZ  sky130_fd_pr__res_xhigh_po_0p35_PYW3KZ_0
timestamp 1716692466
transform 0 1 14202 -1 0 39763
box -201 -4582 201 4582
use sky130_fd_pr__res_xhigh_po_0p35_QMT3WJ  sky130_fd_pr__res_xhigh_po_0p35_QMT3WJ_0
timestamp 1717301720
transform 0 1 5142 -1 0 39763
box -201 -4582 201 4582
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1707688321
transform 1 0 3128 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_17
timestamp 1707688321
transform 1 0 5704 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_18
timestamp 1707688321
transform 1 0 8280 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_19
timestamp 1707688321
transform 1 0 10856 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_20
timestamp 1707688321
transform 1 0 13432 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_21
timestamp 1707688321
transform 1 0 16008 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_22
timestamp 1707688321
transform 1 0 18584 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_23
timestamp 1707688321
transform 1 0 21160 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_24
timestamp 1707688321
transform 1 0 23736 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_25
timestamp 1707688321
transform 1 0 26312 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 1707688321
transform 1 0 28888 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_27
timestamp 1707688321
transform 1 0 5704 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp 1707688321
transform 1 0 10856 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_29
timestamp 1707688321
transform 1 0 16008 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 1707688321
transform 1 0 21160 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_31
timestamp 1707688321
transform 1 0 26312 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_32
timestamp 1707688321
transform 1 0 3128 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_33
timestamp 1707688321
transform 1 0 8280 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_34
timestamp 1707688321
transform 1 0 13432 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_35
timestamp 1707688321
transform 1 0 18584 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_36
timestamp 1707688321
transform 1 0 23736 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_37
timestamp 1707688321
transform 1 0 28888 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_38
timestamp 1707688321
transform 1 0 5704 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_39
timestamp 1707688321
transform 1 0 10856 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1707688321
transform 1 0 16008 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_41
timestamp 1707688321
transform 1 0 21160 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 1707688321
transform 1 0 26312 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp 1707688321
transform 1 0 3128 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_44
timestamp 1707688321
transform 1 0 8280 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_45
timestamp 1707688321
transform 1 0 13432 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_46
timestamp 1707688321
transform 1 0 18584 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_47
timestamp 1707688321
transform 1 0 23736 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_48
timestamp 1707688321
transform 1 0 28888 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_49
timestamp 1707688321
transform 1 0 5704 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_50
timestamp 1707688321
transform 1 0 10856 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_51
timestamp 1707688321
transform 1 0 16008 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_52
timestamp 1707688321
transform 1 0 21160 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_53
timestamp 1707688321
transform 1 0 26312 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_54
timestamp 1707688321
transform 1 0 3128 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 1707688321
transform 1 0 8280 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 1707688321
transform 1 0 13432 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1707688321
transform 1 0 18584 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_58
timestamp 1707688321
transform 1 0 23736 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_59
timestamp 1707688321
transform 1 0 28888 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_60
timestamp 1707688321
transform 1 0 3128 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_61
timestamp 1707688321
transform 1 0 5704 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp 1707688321
transform 1 0 8280 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp 1707688321
transform 1 0 10856 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_64
timestamp 1707688321
transform 1 0 13432 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_65
timestamp 1707688321
transform 1 0 16008 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_66
timestamp 1707688321
transform 1 0 18584 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_67
timestamp 1707688321
transform 1 0 21160 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_68
timestamp 1707688321
transform 1 0 23736 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_69
timestamp 1707688321
transform 1 0 26312 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_70
timestamp 1707688321
transform 1 0 28888 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_9
timestamp 1707688321
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_10
timestamp 1707688321
transform 1 0 5244 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_11
timestamp 1707688321
transform 1 0 4508 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_12
timestamp 1707688321
transform 1 0 3772 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_13
timestamp 1707688321
transform 1 0 3220 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_14
timestamp 1707688321
transform 1 0 2300 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_15
timestamp 1707688321
transform 1 0 1564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_dlmiles_schmitt_playground_16
timestamp 1707688321
transform 1 0 828 0 -1 44608
box -38 -48 314 592
<< labels >>
flabel metal4 15940 40208 16260 44656 0 FreeSans 1920 90 0 0 VGND
flabel metal4 23714 40208 24034 44656 0 FreeSans 1920 90 0 0 VGND
flabel metal4 4279 40208 4599 44656 0 FreeSans 1920 90 0 0 VPWR
flabel metal4 12053 40208 12373 44656 0 FreeSans 1920 90 0 0 VPWR
flabel metal4 27601 40208 27921 44656 0 FreeSans 1920 90 0 0 VPWR
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 28766 39604 28826 39804 0 FreeSans 480 90 0 0 oa_ctrl[0]
port 4 nsew signal tristate
flabel metal4 s 12574 39604 12634 39804 0 FreeSans 480 90 0 0 oa_ctrl[10]
port 5 nsew signal tristate
flabel metal4 s 9630 39604 9690 39804 0 FreeSans 480 90 0 0 oa_ctrl[12]
port 7 nsew signal tristate
flabel metal4 s 7273 39604 7333 39804 0 FreeSans 480 90 0 0 oa_ctrl[13]
port 8 nsew signal tristate
flabel metal4 s 5801 39604 5861 39804 0 FreeSans 480 90 0 0 oa_ctrl[14]
port 9 nsew signal tristate
flabel metal4 s 4329 39604 4389 39804 0 FreeSans 480 90 0 0 oa_ctrl[15]
port 10 nsew signal tristate
flabel metal4 s 27294 39604 27354 39804 0 FreeSans 480 90 0 0 oa_ctrl[1]
port 11 nsew signal tristate
flabel metal4 s 25822 39604 25882 39804 0 FreeSans 480 90 0 0 oa_ctrl[2]
port 12 nsew signal tristate
flabel metal4 s 24350 39604 24410 39804 0 FreeSans 480 90 0 0 oa_ctrl[3]
port 13 nsew signal tristate
flabel metal4 s 22878 39604 22938 39804 0 FreeSans 480 90 0 0 oa_ctrl[4]
port 14 nsew signal tristate
flabel metal4 s 21406 39604 21466 39804 0 FreeSans 480 90 0 0 oa_ctrl[5]
port 15 nsew signal tristate
flabel metal4 s 18462 39604 18522 39804 0 FreeSans 480 90 0 0 oa_ctrl[6]
port 16 nsew signal tristate
flabel metal4 s 16990 39604 17050 39804 0 FreeSans 480 90 0 0 oa_ctrl[7]
port 17 nsew signal tristate
flabel metal4 s 15518 39604 15578 39804 0 FreeSans 480 90 0 0 oa_ctrl[8]
port 18 nsew signal tristate
flabel metal4 s 14046 39604 14106 39804 0 FreeSans 480 90 0 0 oa_ctrl[9]
port 19 nsew signal tristate
flabel metal4 s 30238 39604 30298 39804 0 FreeSans 480 90 0 0 oa_ena
port 20 nsew signal tristate
flabel metal4 s 2857 39604 2917 39804 0 FreeSans 480 90 0 0 oa_por[0]
port 21 nsew signal tristate
flabel metal4 s 1385 39604 1445 39804 0 FreeSans 480 90 0 0 oa_por[1]
port 22 nsew signal tristate
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 23 nsew signal input
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 24 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 25 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 26 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 27 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 28 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 29 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 30 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 31 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 32 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 33 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 34 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 35 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 36 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 37 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 38 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 39 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 40 nsew signal tristate
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 41 nsew signal tristate
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 42 nsew signal tristate
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 43 nsew signal tristate
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 44 nsew signal tristate
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 45 nsew signal tristate
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 46 nsew signal tristate
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 47 nsew signal tristate
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 48 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 49 nsew signal tristate
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 50 nsew signal tristate
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 51 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 52 nsew signal tristate
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 53 nsew signal tristate
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 54 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 55 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 56 nsew signal tristate
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 57 nsew signal tristate
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 58 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 59 nsew signal tristate
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 60 nsew signal tristate
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 61 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 62 nsew signal tristate
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 63 nsew signal tristate
flabel metal4 200 1000 520 44152 0 FreeSans 1440 90 0 0 VPWR
port 64 nsew power bidirectional
flabel metal4 31488 1000 31808 44656 0 FreeSans 1440 90 0 0 VGND
port 65 nsew ground bidirectional
flabel metal4 31282 0 31462 200 0 FreeSans 400 0 0 0 ua[0]
port 66 nsew signal bidirectional
flabel metal4 26866 0 27046 200 0 FreeSans 400 0 0 0 ua[1]
port 67 nsew signal bidirectional
flabel metal4 22450 0 22630 200 0 FreeSans 400 0 0 0 ua[2]
port 68 nsew signal bidirectional
flabel metal4 18034 0 18214 200 0 FreeSans 400 0 0 0 ua[3]
port 69 nsew signal bidirectional
flabel metal4 13618 0 13798 200 0 FreeSans 400 0 0 0 ua[4]
port 70 nsew signal bidirectional
flabel metal4 9202 0 9382 200 0 FreeSans 400 0 0 0 ua[5]
port 71 nsew signal bidirectional
flabel metal4 4786 0 4966 200 0 FreeSans 400 0 0 0 ua[6]
port 72 nsew signal bidirectional
flabel metal4 370 0 550 200 0 FreeSans 400 0 0 0 ua[7]
port 73 nsew signal bidirectional
flabel metal4 s 11102 39604 11162 39804 0 FreeSans 480 90 0 0 oa_ctrl[11]
port 6 nsew signal tristate
flabel metal4 19827 1000 20147 44656 0 FreeSans 1440 90 0 0 VPWR
port 64 nsew power bidirectional
flabel metal4 8166 1000 8486 44656 0 FreeSans 1440 90 0 0 VGND
port 65 nsew ground bidirectional
flabel metal2 4342 41062 4528 41114 0 FreeSans 400 0 0 0 patch_por0
flabel metal2 2134 41062 2320 41114 0 FreeSans 400 0 0 0 patch_por1
flabel space 21000 41922 21130 42171 0 FreeSans 400 0 0 0 patch_filler_0_3_222
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
