magic
tech sky130A
magscale 1 2
timestamp 1717291860
<< metal3 >>
rect 26856 1030 30238 1040
rect 26856 850 26870 1030
rect 27045 850 30050 1030
rect 30230 850 30240 1030
rect 26856 840 30238 850
rect 24690 630 24890 640
rect 24690 450 24700 630
rect 24880 450 24890 630
rect 24690 440 24890 450
rect 24690 430 31472 440
rect 24690 250 31280 430
rect 31460 250 31472 430
rect 24690 240 31472 250
<< via3 >>
rect 26870 850 27045 1030
rect 30050 850 30230 1030
rect 24700 450 24880 630
rect 31280 250 31460 430
<< metal4 >>
rect 1770 640 1970 1200
rect 26856 1030 27056 1040
rect 26856 850 26870 1030
rect 27045 850 27056 1030
rect 1770 630 24890 640
rect 1770 450 24700 630
rect 24880 450 24890 630
rect 1770 440 24890 450
rect 26856 0 27056 850
rect 30038 1030 30238 1198
rect 30038 850 30050 1030
rect 30230 850 30238 1030
rect 30038 840 30238 850
rect 31272 430 31472 440
rect 31272 250 31280 430
rect 31460 250 31472 430
rect 31272 0 31472 250
<< properties >>
string FIXED_BBOX 0 0 32200 1200
<< end >>
