//
//

`ifdef SYNTHESIS

`define TT_ANALOG_POWER 1

`define TT_ANALOG_INTERNAL_SIGNAL_PORTS 1

`endif
