magic
tech sky130A
magscale 1 2
timestamp 1717261669
<< locali >>
rect 0 2085 1950 2100
rect 0 492 43 2085
rect 87 2033 1950 2085
rect 87 532 170 2033
rect 300 532 1490 533
rect 87 492 1490 532
rect 0 294 15 492
rect 1427 294 1490 492
rect 0 68 1490 294
rect 1775 68 1950 2033
rect 0 0 1950 68
rect 1985 2086 3673 2100
rect 1985 1612 3163 2086
rect 1985 73 2160 1612
rect 2998 533 3163 1612
rect 2445 489 3163 533
rect 3207 489 3673 2086
rect 2445 294 2653 489
rect 3657 294 3673 489
rect 2445 73 3673 294
rect 1985 0 3673 73
<< viali >>
rect 43 492 87 2085
rect 15 294 1427 492
rect 3163 489 3207 2086
rect 2653 294 3657 489
<< metal1 >>
rect 30 2085 100 2097
rect 30 499 43 2085
rect 3 492 43 499
rect 87 499 100 2085
rect 3150 2086 3220 2097
rect 130 1981 200 1987
rect 130 1923 136 1981
rect 194 1977 200 1981
rect 194 1923 1920 1977
rect 130 1917 1920 1923
rect 245 1432 287 1873
rect 235 1152 245 1432
rect 317 1152 327 1432
rect 245 689 287 1152
rect 373 992 415 1873
rect 501 1432 543 1873
rect 490 1152 500 1432
rect 572 1152 582 1432
rect 365 712 375 992
rect 447 712 457 992
rect 373 689 415 712
rect 501 689 543 1152
rect 629 992 671 1873
rect 757 1432 799 1873
rect 745 1152 755 1432
rect 827 1152 837 1432
rect 623 712 633 992
rect 705 712 715 992
rect 629 689 671 712
rect 757 689 799 1152
rect 885 992 927 1873
rect 1013 1432 1055 1873
rect 1000 1152 1010 1432
rect 1082 1152 1092 1432
rect 878 712 888 992
rect 960 712 970 992
rect 885 689 927 712
rect 1013 689 1055 1152
rect 1141 992 1183 1873
rect 1269 1432 1311 1873
rect 1255 1152 1265 1432
rect 1337 1152 1347 1432
rect 1133 712 1143 992
rect 1215 712 1225 992
rect 1141 689 1183 712
rect 1269 689 1311 1152
rect 1397 992 1439 1873
rect 1525 1432 1567 1873
rect 1510 1152 1520 1432
rect 1592 1152 1602 1432
rect 1388 712 1398 992
rect 1470 712 1480 992
rect 1397 689 1439 712
rect 1525 689 1567 1152
rect 1653 992 1695 1873
rect 1643 712 1653 992
rect 1725 712 1735 992
rect 1653 689 1695 712
rect 1840 642 1920 1917
rect 2290 1502 3120 1562
rect 2238 1432 2280 1462
rect 2225 1152 2235 1432
rect 2307 1152 2317 1432
rect 2238 682 2280 1152
rect 2366 992 2408 1462
rect 2494 1432 2536 1462
rect 2480 1152 2490 1432
rect 2562 1152 2572 1432
rect 2358 712 2368 992
rect 2440 712 2450 992
rect 2366 682 2408 712
rect 2494 682 2536 1152
rect 2622 992 2664 1462
rect 2750 1432 2792 1462
rect 2735 1152 2745 1432
rect 2817 1152 2827 1432
rect 2613 712 2623 992
rect 2695 712 2705 992
rect 2622 682 2664 712
rect 2750 682 2792 1152
rect 2878 992 2920 1462
rect 2870 712 2880 992
rect 2932 712 2942 992
rect 2878 682 2920 712
rect 3066 642 3120 1502
rect 300 582 1920 642
rect 2290 582 3120 642
rect 87 492 1440 499
rect 3 294 8 492
rect 1427 294 1440 492
rect 1567 402 1607 411
rect 1655 402 1695 411
rect 1840 402 1920 582
rect 2239 402 2279 405
rect 2327 402 2367 405
rect 1543 332 1553 402
rect 1605 332 1615 402
rect 1648 332 1658 402
rect 1710 332 1720 402
rect 1830 332 1840 402
rect 1920 332 1930 402
rect 2213 332 2223 402
rect 2275 332 2285 402
rect 2318 332 2328 402
rect 2380 332 2390 402
rect 3 286 1440 294
rect 1567 229 1607 332
rect 1655 229 1695 332
rect 1840 322 1920 332
rect 2239 223 2279 332
rect 2327 223 2367 332
rect 2550 193 2610 582
rect 3150 499 3163 2086
rect 2640 492 3163 499
rect 3207 499 3220 2086
rect 3207 492 3670 499
rect 2640 489 3028 492
rect 3232 489 3670 492
rect 2640 484 2653 489
rect 2640 342 2650 484
rect 2640 294 2653 342
rect 3659 335 3670 489
rect 3657 294 3670 335
rect 2640 292 3028 294
rect 3232 292 3670 294
rect 2640 286 3670 292
rect 1210 184 1290 192
rect 1210 130 1218 184
rect 1282 182 1290 184
rect 2539 187 2621 193
rect 2539 182 2545 187
rect 1282 132 2545 182
rect 1282 130 1290 132
rect 1210 122 1290 130
rect 2539 127 2545 132
rect 2615 127 2621 187
rect 2539 121 2621 127
<< via1 >>
rect 136 1923 194 1981
rect 245 1152 317 1432
rect 500 1152 572 1432
rect 375 712 447 992
rect 755 1152 827 1432
rect 633 712 705 992
rect 1010 1152 1082 1432
rect 888 712 960 992
rect 1265 1152 1337 1432
rect 1143 712 1215 992
rect 1520 1152 1592 1432
rect 1398 712 1470 992
rect 1653 712 1725 992
rect 2235 1152 2307 1432
rect 2490 1152 2562 1432
rect 2368 712 2440 992
rect 2745 1152 2817 1432
rect 2623 712 2695 992
rect 2880 712 2932 992
rect 8 294 15 492
rect 15 294 192 492
rect 1343 342 1427 482
rect 1553 332 1605 402
rect 1658 332 1710 402
rect 1840 332 1920 402
rect 2223 332 2275 402
rect 2328 332 2380 402
rect 3028 489 3163 492
rect 3163 489 3207 492
rect 3207 489 3232 492
rect 2650 342 2653 484
rect 2653 342 2730 484
rect 3028 294 3232 489
rect 3588 335 3657 489
rect 3657 335 3659 489
rect 3028 292 3232 294
rect 1218 130 1282 184
rect 2545 127 2615 187
<< metal2 >>
rect 0 1981 200 2002
rect 0 1923 136 1981
rect 194 1923 200 1981
rect 0 1802 200 1923
rect 0 1432 2817 1442
rect 0 1152 245 1432
rect 317 1152 500 1432
rect 572 1152 755 1432
rect 827 1152 1010 1432
rect 1082 1152 1265 1432
rect 1337 1152 1520 1432
rect 1592 1152 2235 1432
rect 2307 1152 2490 1432
rect 2562 1152 2745 1432
rect 0 1142 2817 1152
rect 370 993 3510 1002
rect 370 992 3319 993
rect 0 682 210 902
rect 370 712 375 992
rect 447 712 633 992
rect 705 712 888 992
rect 960 712 1143 992
rect 1215 712 1398 992
rect 1470 712 1653 992
rect 1725 712 2368 992
rect 2440 712 2623 992
rect 2695 712 2880 992
rect 2932 712 3319 992
rect 370 711 3319 712
rect 3501 711 3510 993
rect 370 702 3510 711
rect 150 602 210 682
rect 150 542 380 602
rect 0 492 210 502
rect 0 294 8 492
rect 192 294 210 492
rect 320 362 380 542
rect 1343 482 1427 492
rect 320 302 1280 362
rect 2640 484 2740 494
rect 1553 402 1605 412
rect 1658 402 1710 412
rect 1840 402 1920 412
rect 2223 402 2275 412
rect 2328 402 2380 412
rect 2640 402 2650 484
rect 1427 342 1553 402
rect 1343 332 1553 342
rect 1650 332 1658 402
rect 1710 332 1840 402
rect 1920 332 2223 402
rect 2275 332 2280 402
rect 2325 332 2328 402
rect 2380 342 2650 402
rect 2730 342 2740 484
rect 2380 332 2740 342
rect 3020 492 3240 500
rect 1553 322 1605 332
rect 1658 322 1710 332
rect 1840 322 1920 332
rect 2223 322 2275 332
rect 2328 322 2380 332
rect 0 282 210 294
rect 1220 192 1280 302
rect 3020 292 3028 492
rect 3232 292 3240 492
rect 3580 489 3667 497
rect 3580 335 3588 489
rect 3659 335 3667 489
rect 3580 327 3667 335
rect 3020 284 3240 292
rect 4193 197 4226 2100
rect 1210 184 1290 192
rect 1210 130 1218 184
rect 1282 130 1290 184
rect 1210 122 1290 130
rect 2536 187 2624 196
rect 2536 127 2545 187
rect 2615 127 2624 187
rect 2536 118 2624 127
rect 4150 187 4226 197
rect 4150 127 4156 187
rect 4220 127 4226 187
rect 4150 117 4226 127
rect 4258 0 4291 2100
rect 4323 0 4356 2100
rect 4388 0 4421 2100
rect 4453 0 4486 2100
rect 4518 0 4551 2100
rect 4583 0 4616 2100
rect 4648 0 4681 2100
rect 4713 0 4746 2100
<< via2 >>
rect 3319 711 3501 993
rect 3036 295 3230 489
rect 3590 337 3657 487
rect 2545 127 2615 187
rect 4156 127 4220 187
<< metal3 >>
rect 3310 993 3510 1012
rect 3310 711 3319 993
rect 3501 711 3510 993
rect 3310 692 3510 711
rect 3025 489 5080 497
rect 3025 295 3033 489
rect 3238 487 4788 489
rect 3238 482 3590 487
rect 3238 342 3582 482
rect 3238 337 3590 342
rect 3657 337 4788 487
rect 3238 335 4788 337
rect 5072 335 5080 489
rect 3238 327 5080 335
rect 3238 295 3240 327
rect 3025 287 3240 295
rect 2536 189 2667 196
rect 2536 125 2541 189
rect 2617 125 2667 189
rect 2536 118 2667 125
rect 2730 189 4230 192
rect 2730 125 2740 189
rect 2817 187 4230 189
rect 2817 127 4156 187
rect 4220 127 4230 187
rect 2817 125 4230 127
rect 2730 122 4230 125
<< via3 >>
rect 3320 712 3500 992
rect 3033 295 3036 489
rect 3036 295 3230 489
rect 3230 295 3238 489
rect 3582 342 3590 482
rect 3590 342 3646 482
rect 4788 335 5072 489
rect 2541 187 2617 189
rect 2541 127 2545 187
rect 2545 127 2615 187
rect 2615 127 2617 187
rect 2541 125 2617 127
rect 2740 125 2817 189
<< metal4 >>
rect 3180 497 3240 2100
rect 3025 489 3240 497
rect 3025 295 3033 489
rect 3238 295 3240 489
rect 3025 287 3240 295
rect 2536 189 2822 192
rect 2536 125 2541 189
rect 2617 125 2740 189
rect 2817 125 2822 189
rect 2536 122 2822 125
rect 3180 0 3240 287
rect 3310 992 3510 2100
rect 3310 712 3320 992
rect 3500 712 3510 992
rect 3310 0 3510 712
rect 3580 497 3640 2100
rect 4780 497 5080 2100
rect 3580 489 5080 497
rect 3580 482 4788 489
rect 3580 342 3582 482
rect 3646 342 4788 482
rect 3580 335 4788 342
rect 5072 335 5080 489
rect 3580 327 5080 335
rect 3580 0 3640 327
rect 4780 0 5080 327
use sky130_fd_pr__nfet_01v8_9BJ5NV#07tgo  sky130_fd_pr__nfet_01v8_9BJ5NV_0_07tgo
timestamp 1716692466
transform 1 0 2303 0 1 283
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_X62NDW#07tgo  sky130_fd_pr__nfet_01v8_lvt_X62NDW_0_07tgo
timestamp 1716692466
transform 1 0 2579 0 1 1072
box -487 -610 487 610
use sky130_fd_pr__pfet_01v8_L75DJ9#07tgo  sky130_fd_pr__pfet_01v8_L75DJ9_0_07tgo
timestamp 1717177448
transform 1 0 1631 0 1 284
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_lvt_E3P74E#07tgo  sky130_fd_pr__pfet_01v8_lvt_E3P74E_0_07tgo
timestamp 1716692466
transform 1 0 971 0 1 1281
box -871 -819 871 819
<< labels >>
flabel metal2 0 692 200 892 0 FreeSans 400 0 0 0 EN
port 6 nsew signal output
flabel metal2 0 1802 200 2002 0 FreeSans 400 0 0 0 EN_N
port 5 nsew signal output
flabel metal2 0 293 200 493 0 FreeSans 400 0 0 0 VPWR
port 2 nsew power bidirectional
flabel via1 3030 292 3230 492 0 FreeSans 400 0 0 0 VGND
port 1 nsew power bidirectional
flabel metal4 4780 327 5080 497 0 FreeSans 400 0 0 0 VGND
port 1 nsew power bidirectional
flabel metal2 3310 702 3510 1002 0 FreeSans 400 0 0 0 AOUT
port 3 nsew signal output
flabel metal2 0 1142 200 1442 0 FreeSans 400 0 0 0 AIN
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 5080 2100
<< end >>
