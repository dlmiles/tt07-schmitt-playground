VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_dlmiles_schmitt_playground
  CLASS BLOCK ;
  FOREIGN tt_um_dlmiles_schmitt_playground ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.600 220.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.135 5.000 100.735 223.280 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 157.440 5.000 159.040 223.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.830 5.000 42.430 223.280 ;
    END
  END VGND
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 222.720001 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 222.720001 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  OBS
      LAYER pwell ;
        RECT 2.905 222.935 3.075 223.125 ;
        RECT 4.285 222.955 4.455 223.125 ;
        RECT 5.665 222.935 5.835 223.125 ;
        RECT 7.500 222.985 7.620 223.095 ;
        RECT 7.965 222.955 8.135 223.125 ;
        RECT 9.345 222.935 9.515 223.125 ;
        RECT 11.180 222.985 11.300 223.095 ;
        RECT 11.645 222.955 11.815 223.125 ;
        RECT 13.025 222.935 13.195 223.125 ;
        RECT 16.245 222.955 16.415 223.125 ;
        RECT 17.625 222.935 17.795 223.125 ;
        RECT 19.005 222.955 19.175 223.125 ;
        RECT 20.385 222.935 20.555 223.125 ;
        RECT 22.220 222.985 22.340 223.095 ;
        RECT 22.685 222.955 22.855 223.125 ;
        RECT 24.065 222.935 24.235 223.125 ;
        RECT 25.900 222.985 26.020 223.095 ;
        RECT 26.365 222.955 26.535 223.125 ;
        RECT 27.755 222.980 27.915 223.090 ;
        RECT 29.135 222.980 29.295 223.090 ;
        RECT 30.045 222.955 30.215 223.125 ;
        RECT 31.425 222.935 31.595 223.125 ;
        RECT 36.945 222.935 37.115 223.125 ;
        RECT 40.635 222.980 40.795 223.090 ;
        RECT 42.005 222.935 42.175 223.125 ;
        RECT 47.525 222.935 47.695 223.125 ;
        RECT 53.045 222.935 53.215 223.125 ;
        RECT 54.885 222.935 55.055 223.125 ;
        RECT 57.640 222.985 57.760 223.095 ;
        RECT 61.780 222.935 61.950 223.125 ;
        RECT 62.240 222.985 62.360 223.095 ;
        RECT 65.925 222.935 66.095 223.125 ;
        RECT 66.395 222.980 66.555 223.090 ;
        RECT 69.600 222.935 69.770 223.125 ;
        RECT 71.445 222.935 71.615 223.125 ;
        RECT 71.905 222.935 72.075 223.125 ;
        RECT 79.725 222.935 79.895 223.125 ;
        RECT 80.655 222.980 80.815 223.090 ;
        RECT 81.570 222.935 81.740 223.125 ;
        RECT 85.705 222.935 85.875 223.125 ;
        RECT 87.085 222.935 87.255 223.125 ;
        RECT 90.765 222.935 90.935 223.125 ;
        RECT 92.600 222.985 92.720 223.095 ;
        RECT 93.525 222.935 93.695 223.125 ;
        RECT 96.285 222.935 96.455 223.125 ;
        RECT 97.665 222.935 97.835 223.125 ;
        RECT 103.185 222.935 103.355 223.125 ;
        RECT 109.625 222.935 109.795 223.125 ;
        RECT 110.085 222.935 110.255 223.125 ;
        RECT 111.465 222.935 111.635 223.125 ;
        RECT 113.300 222.985 113.420 223.095 ;
        RECT 113.765 222.955 113.935 223.125 ;
        RECT 113.765 222.935 113.965 222.955 ;
        RECT 117.445 222.935 117.615 223.125 ;
        RECT 119.285 222.935 119.455 223.125 ;
        RECT 122.965 222.955 123.135 223.125 ;
        RECT 122.985 222.935 123.135 222.955 ;
        RECT 126.185 222.935 126.355 223.125 ;
        RECT 127.565 222.935 127.735 223.125 ;
        RECT 128.025 222.935 128.195 223.125 ;
        RECT 132.175 222.980 132.335 223.090 ;
        RECT 134.005 222.935 134.175 223.125 ;
        RECT 134.740 222.935 134.910 223.125 ;
        RECT 141.825 222.935 141.995 223.125 ;
        RECT 143.205 222.935 143.375 223.125 ;
        RECT 143.675 222.980 143.835 223.090 ;
        RECT 148.450 222.935 148.620 223.125 ;
        RECT 152.590 222.935 152.760 223.125 ;
        RECT 156.545 222.935 156.715 223.125 ;
        RECT 157.925 222.935 158.095 223.125 ;
        RECT 2.765 222.125 4.135 222.935 ;
        RECT 5.525 222.125 7.355 222.935 ;
        RECT 9.205 222.125 11.035 222.935 ;
        RECT 12.885 222.125 15.635 222.935 ;
        RECT 15.655 222.065 16.085 222.850 ;
        RECT 17.485 222.125 18.855 222.935 ;
        RECT 20.245 222.125 22.075 222.935 ;
        RECT 23.925 222.125 25.755 222.935 ;
        RECT 28.535 222.065 28.965 222.850 ;
        RECT 31.285 222.125 36.795 222.935 ;
        RECT 36.805 222.125 40.475 222.935 ;
        RECT 41.415 222.065 41.845 222.850 ;
        RECT 41.865 222.125 47.375 222.935 ;
        RECT 47.385 222.125 52.895 222.935 ;
        RECT 52.905 222.125 54.275 222.935 ;
        RECT 54.295 222.065 54.725 222.850 ;
        RECT 54.745 222.125 57.495 222.935 ;
        RECT 58.205 222.025 62.095 222.935 ;
        RECT 62.565 222.255 66.235 222.935 ;
        RECT 62.565 222.025 63.495 222.255 ;
        RECT 67.175 222.065 67.605 222.850 ;
        RECT 67.725 222.025 69.915 222.935 ;
        RECT 69.925 222.255 71.755 222.935 ;
        RECT 69.925 222.025 71.270 222.255 ;
        RECT 71.765 222.125 77.275 222.935 ;
        RECT 77.295 222.025 80.025 222.935 ;
        RECT 80.055 222.065 80.485 222.850 ;
        RECT 81.425 222.025 85.315 222.935 ;
        RECT 85.565 222.125 86.935 222.935 ;
        RECT 87.055 222.255 90.520 222.935 ;
        RECT 89.600 222.025 90.520 222.255 ;
        RECT 90.625 222.125 92.455 222.935 ;
        RECT 92.935 222.065 93.365 222.850 ;
        RECT 93.395 222.025 96.125 222.935 ;
        RECT 96.155 222.025 97.505 222.935 ;
        RECT 97.525 222.125 103.035 222.935 ;
        RECT 103.045 222.125 105.795 222.935 ;
        RECT 105.815 222.065 106.245 222.850 ;
        RECT 106.360 222.255 109.825 222.935 ;
        RECT 106.360 222.025 107.280 222.255 ;
        RECT 109.955 222.025 111.305 222.935 ;
        RECT 111.325 222.125 113.155 222.935 ;
        RECT 113.765 222.255 117.295 222.935 ;
        RECT 114.470 222.025 117.295 222.255 ;
        RECT 117.305 222.125 118.675 222.935 ;
        RECT 118.695 222.065 119.125 222.850 ;
        RECT 119.145 222.125 122.815 222.935 ;
        RECT 122.985 222.115 124.915 222.935 ;
        RECT 125.125 222.155 126.495 222.935 ;
        RECT 126.505 222.155 127.875 222.935 ;
        RECT 127.885 222.125 131.555 222.935 ;
        RECT 123.965 222.025 124.915 222.115 ;
        RECT 131.575 222.065 132.005 222.850 ;
        RECT 132.945 222.155 134.315 222.935 ;
        RECT 134.325 222.255 138.225 222.935 ;
        RECT 138.560 222.255 142.025 222.935 ;
        RECT 134.325 222.025 135.255 222.255 ;
        RECT 138.560 222.025 139.480 222.255 ;
        RECT 142.145 222.155 143.515 222.935 ;
        RECT 144.455 222.065 144.885 222.850 ;
        RECT 145.135 222.255 149.035 222.935 ;
        RECT 149.275 222.255 153.175 222.935 ;
        RECT 148.105 222.025 149.035 222.255 ;
        RECT 152.245 222.025 153.175 222.255 ;
        RECT 153.280 222.255 156.745 222.935 ;
        RECT 153.280 222.025 154.200 222.255 ;
        RECT 156.865 222.125 158.235 222.935 ;
      LAYER nwell ;
        RECT 2.570 218.905 158.430 221.735 ;
      LAYER pwell ;
        RECT 2.765 217.705 4.135 218.515 ;
        RECT 4.145 217.705 9.655 218.515 ;
        RECT 9.665 217.705 15.175 218.515 ;
        RECT 15.655 217.790 16.085 218.575 ;
        RECT 16.105 217.705 21.615 218.515 ;
        RECT 21.625 217.705 27.135 218.515 ;
        RECT 27.145 217.705 32.655 218.515 ;
        RECT 32.665 217.705 38.175 218.515 ;
        RECT 38.185 217.705 40.935 218.515 ;
        RECT 41.415 217.790 41.845 218.575 ;
        RECT 41.865 217.705 47.375 218.515 ;
        RECT 47.385 217.705 52.895 218.515 ;
        RECT 52.905 217.705 54.275 218.515 ;
        RECT 54.295 217.705 55.645 218.615 ;
        RECT 61.940 218.385 62.850 218.605 ;
        RECT 64.385 218.385 65.735 218.615 ;
        RECT 55.675 217.705 58.415 218.385 ;
        RECT 58.425 217.705 65.735 218.385 ;
        RECT 65.785 217.705 67.155 218.515 ;
        RECT 67.175 217.790 67.605 218.575 ;
        RECT 67.635 217.705 70.375 218.385 ;
        RECT 70.625 217.705 74.515 218.615 ;
        RECT 74.995 217.705 76.345 218.615 ;
        RECT 76.375 217.705 79.105 218.615 ;
        RECT 82.640 218.385 83.550 218.605 ;
        RECT 85.085 218.385 86.855 218.615 ;
        RECT 79.125 217.705 86.855 218.385 ;
        RECT 87.185 217.705 91.075 218.615 ;
        RECT 91.085 217.705 92.915 218.515 ;
        RECT 92.935 217.790 93.365 218.575 ;
        RECT 96.040 218.385 96.960 218.615 ;
        RECT 93.495 217.705 96.960 218.385 ;
        RECT 97.075 217.705 99.805 218.615 ;
        RECT 103.800 218.385 104.710 218.605 ;
        RECT 106.245 218.385 107.595 218.615 ;
        RECT 100.285 217.705 107.595 218.385 ;
        RECT 107.685 218.385 109.035 218.615 ;
        RECT 110.570 218.385 111.480 218.605 ;
        RECT 115.850 218.385 118.675 218.615 ;
        RECT 107.685 217.705 114.995 218.385 ;
        RECT 115.145 217.705 118.675 218.385 ;
        RECT 118.695 217.790 119.125 218.575 ;
        RECT 119.155 217.705 120.505 218.615 ;
        RECT 124.960 218.385 125.870 218.605 ;
        RECT 127.405 218.385 128.755 218.615 ;
        RECT 121.445 217.705 128.755 218.385 ;
        RECT 128.805 217.705 132.475 218.515 ;
        RECT 136.460 218.385 137.370 218.605 ;
        RECT 138.905 218.385 140.255 218.615 ;
        RECT 143.505 218.385 144.435 218.615 ;
        RECT 132.945 217.705 140.255 218.385 ;
        RECT 140.535 217.705 144.435 218.385 ;
        RECT 144.455 217.790 144.885 218.575 ;
        RECT 148.420 218.385 149.330 218.605 ;
        RECT 150.865 218.385 152.215 218.615 ;
        RECT 144.905 217.705 152.215 218.385 ;
        RECT 152.820 218.385 153.740 218.615 ;
        RECT 152.820 217.705 156.285 218.385 ;
        RECT 156.865 217.705 158.235 218.515 ;
        RECT 2.905 217.495 3.075 217.705 ;
        RECT 4.285 217.495 4.455 217.705 ;
        RECT 9.805 217.495 9.975 217.705 ;
        RECT 15.325 217.655 15.495 217.685 ;
        RECT 15.320 217.545 15.495 217.655 ;
        RECT 15.325 217.495 15.495 217.545 ;
        RECT 16.245 217.515 16.415 217.705 ;
        RECT 20.845 217.495 21.015 217.685 ;
        RECT 21.765 217.515 21.935 217.705 ;
        RECT 26.365 217.495 26.535 217.685 ;
        RECT 27.285 217.515 27.455 217.705 ;
        RECT 28.200 217.545 28.320 217.655 ;
        RECT 29.125 217.495 29.295 217.685 ;
        RECT 32.805 217.515 32.975 217.705 ;
        RECT 34.645 217.495 34.815 217.685 ;
        RECT 38.325 217.515 38.495 217.705 ;
        RECT 40.165 217.495 40.335 217.685 ;
        RECT 41.080 217.545 41.200 217.655 ;
        RECT 42.005 217.515 42.175 217.705 ;
        RECT 45.685 217.495 45.855 217.685 ;
        RECT 47.525 217.515 47.695 217.705 ;
        RECT 51.205 217.495 51.375 217.685 ;
        RECT 53.045 217.515 53.215 217.705 ;
        RECT 53.960 217.545 54.080 217.655 ;
        RECT 54.425 217.515 54.595 217.705 ;
        RECT 54.885 217.495 55.055 217.685 ;
        RECT 58.105 217.515 58.275 217.705 ;
        RECT 58.565 217.515 58.735 217.705 ;
        RECT 65.465 217.495 65.635 217.685 ;
        RECT 65.925 217.495 66.095 217.705 ;
        RECT 70.065 217.515 70.235 217.705 ;
        RECT 74.200 217.685 74.370 217.705 ;
        RECT 74.200 217.515 74.375 217.685 ;
        RECT 74.665 217.655 74.835 217.685 ;
        RECT 74.660 217.545 74.835 217.655 ;
        RECT 74.665 217.515 74.835 217.545 ;
        RECT 75.125 217.515 75.295 217.705 ;
        RECT 76.505 217.515 76.675 217.705 ;
        RECT 77.895 217.540 78.055 217.650 ;
        RECT 74.205 217.495 74.375 217.515 ;
        RECT 78.805 217.495 78.975 217.685 ;
        RECT 79.265 217.515 79.435 217.705 ;
        RECT 80.645 217.495 80.815 217.685 ;
        RECT 90.760 217.515 90.930 217.705 ;
        RECT 91.225 217.515 91.395 217.705 ;
        RECT 93.525 217.515 93.695 217.705 ;
        RECT 95.365 217.495 95.535 217.685 ;
        RECT 95.835 217.540 95.995 217.650 ;
        RECT 96.745 217.495 96.915 217.685 ;
        RECT 97.205 217.515 97.375 217.705 ;
        RECT 99.960 217.545 100.080 217.655 ;
        RECT 100.425 217.515 100.595 217.705 ;
        RECT 106.415 217.540 106.575 217.650 ;
        RECT 107.325 217.495 107.495 217.685 ;
        RECT 114.685 217.515 114.855 217.705 ;
        RECT 115.145 217.685 115.345 217.705 ;
        RECT 115.145 217.515 115.315 217.685 ;
        RECT 116.525 217.495 116.695 217.685 ;
        RECT 117.905 217.495 118.075 217.685 ;
        RECT 120.205 217.515 120.375 217.705 ;
        RECT 120.675 217.550 120.835 217.660 ;
        RECT 121.585 217.515 121.755 217.705 ;
        RECT 126.185 217.495 126.355 217.685 ;
        RECT 126.640 217.545 126.760 217.655 ;
        RECT 127.105 217.495 127.275 217.685 ;
        RECT 128.945 217.515 129.115 217.705 ;
        RECT 132.620 217.545 132.740 217.655 ;
        RECT 133.085 217.495 133.255 217.705 ;
        RECT 133.555 217.540 133.715 217.650 ;
        RECT 135.385 217.495 135.555 217.685 ;
        RECT 135.845 217.495 136.015 217.685 ;
        RECT 143.850 217.515 144.020 217.705 ;
        RECT 144.125 217.495 144.295 217.685 ;
        RECT 145.045 217.515 145.215 217.705 ;
        RECT 145.505 217.495 145.675 217.685 ;
        RECT 146.885 217.495 147.055 217.685 ;
        RECT 147.345 217.495 147.515 217.685 ;
        RECT 152.400 217.545 152.520 217.655 ;
        RECT 155.625 217.495 155.795 217.685 ;
        RECT 156.085 217.515 156.255 217.705 ;
        RECT 156.540 217.545 156.660 217.655 ;
        RECT 157.925 217.495 158.095 217.705 ;
        RECT 2.765 216.685 4.135 217.495 ;
        RECT 4.145 216.685 9.655 217.495 ;
        RECT 9.665 216.685 15.175 217.495 ;
        RECT 15.185 216.685 20.695 217.495 ;
        RECT 20.705 216.685 26.215 217.495 ;
        RECT 26.225 216.685 28.055 217.495 ;
        RECT 28.535 216.625 28.965 217.410 ;
        RECT 28.985 216.685 34.495 217.495 ;
        RECT 34.505 216.685 40.015 217.495 ;
        RECT 40.025 216.685 45.535 217.495 ;
        RECT 45.545 216.685 51.055 217.495 ;
        RECT 51.065 216.685 53.815 217.495 ;
        RECT 54.295 216.625 54.725 217.410 ;
        RECT 54.745 216.685 56.575 217.495 ;
        RECT 56.670 216.815 65.775 217.495 ;
        RECT 65.785 216.815 70.600 217.495 ;
        RECT 70.845 216.815 74.515 217.495 ;
        RECT 74.930 216.815 77.355 217.495 ;
        RECT 70.845 216.585 71.775 216.815 ;
        RECT 78.675 216.585 80.025 217.495 ;
        RECT 80.055 216.625 80.485 217.410 ;
        RECT 80.505 216.815 87.815 217.495 ;
        RECT 84.020 216.595 84.930 216.815 ;
        RECT 86.465 216.585 87.815 216.815 ;
        RECT 87.945 216.815 95.675 217.495 ;
        RECT 96.605 216.815 105.795 217.495 ;
        RECT 87.945 216.585 89.715 216.815 ;
        RECT 91.250 216.595 92.160 216.815 ;
        RECT 101.115 216.595 102.045 216.815 ;
        RECT 104.875 216.585 105.795 216.815 ;
        RECT 105.815 216.625 106.245 217.410 ;
        RECT 107.185 216.815 116.290 217.495 ;
        RECT 116.385 216.685 117.755 217.495 ;
        RECT 117.765 216.815 125.075 217.495 ;
        RECT 121.280 216.595 122.190 216.815 ;
        RECT 123.725 216.585 125.075 216.815 ;
        RECT 125.135 216.585 126.485 217.495 ;
        RECT 126.965 217.265 128.535 217.495 ;
        RECT 130.625 217.455 131.545 217.495 ;
        RECT 130.625 217.265 131.555 217.455 ;
        RECT 126.965 216.905 131.555 217.265 ;
        RECT 126.965 216.815 131.545 216.905 ;
        RECT 128.545 216.585 131.545 216.815 ;
        RECT 131.575 216.625 132.005 217.410 ;
        RECT 132.025 216.715 133.395 217.495 ;
        RECT 134.325 216.715 135.695 217.495 ;
        RECT 135.705 216.685 137.075 217.495 ;
        RECT 137.125 216.815 144.435 217.495 ;
        RECT 137.125 216.585 138.475 216.815 ;
        RECT 140.010 216.595 140.920 216.815 ;
        RECT 144.445 216.715 145.815 217.495 ;
        RECT 145.825 216.715 147.195 217.495 ;
        RECT 147.205 216.815 154.515 217.495 ;
        RECT 150.720 216.595 151.630 216.815 ;
        RECT 153.165 216.585 154.515 216.815 ;
        RECT 154.565 216.715 155.935 217.495 ;
        RECT 156.865 216.685 158.235 217.495 ;
      LAYER nwell ;
        RECT 2.570 213.465 158.430 216.295 ;
      LAYER pwell ;
        RECT 2.765 212.265 4.135 213.075 ;
        RECT 4.145 212.265 9.655 213.075 ;
        RECT 9.665 212.265 15.175 213.075 ;
        RECT 15.655 212.350 16.085 213.135 ;
        RECT 16.105 212.265 21.615 213.075 ;
        RECT 21.625 212.265 27.135 213.075 ;
        RECT 27.145 212.265 32.655 213.075 ;
        RECT 32.665 212.265 38.175 213.075 ;
        RECT 38.185 212.265 40.935 213.075 ;
        RECT 41.415 212.350 41.845 213.135 ;
        RECT 41.865 212.265 47.375 213.075 ;
        RECT 47.385 212.265 52.895 213.075 ;
        RECT 52.905 212.265 54.275 213.075 ;
        RECT 59.815 212.945 62.815 213.175 ;
        RECT 54.295 212.265 57.035 212.945 ;
        RECT 57.055 212.265 59.795 212.945 ;
        RECT 59.815 212.855 64.395 212.945 ;
        RECT 59.805 212.495 64.395 212.855 ;
        RECT 59.805 212.305 60.735 212.495 ;
        RECT 59.815 212.265 60.735 212.305 ;
        RECT 62.825 212.265 64.395 212.495 ;
        RECT 64.405 212.265 67.145 212.945 ;
        RECT 67.175 212.350 67.605 213.135 ;
        RECT 67.865 212.265 71.755 213.175 ;
        RECT 71.765 212.265 73.595 213.075 ;
        RECT 74.090 212.945 77.600 213.175 ;
        RECT 73.605 212.265 77.600 212.945 ;
        RECT 77.985 212.265 81.875 213.175 ;
        RECT 81.970 212.265 91.075 212.945 ;
        RECT 91.085 212.265 92.915 212.945 ;
        RECT 92.935 212.350 93.365 213.135 ;
        RECT 93.385 212.265 98.895 213.075 ;
        RECT 98.905 212.265 101.655 213.075 ;
        RECT 102.125 212.945 103.055 213.175 ;
        RECT 106.360 212.945 107.280 213.175 ;
        RECT 110.040 212.945 110.960 213.175 ;
        RECT 114.470 212.945 117.295 213.175 ;
        RECT 102.125 212.265 106.025 212.945 ;
        RECT 106.360 212.265 109.825 212.945 ;
        RECT 110.040 212.265 113.505 212.945 ;
        RECT 113.765 212.265 117.295 212.945 ;
        RECT 117.305 212.265 118.675 213.045 ;
        RECT 118.695 212.350 119.125 213.135 ;
        RECT 119.145 212.945 120.075 213.175 ;
        RECT 125.420 212.945 126.330 213.165 ;
        RECT 127.865 212.945 129.215 213.175 ;
        RECT 119.145 212.265 121.895 212.945 ;
        RECT 121.905 212.265 129.215 212.945 ;
        RECT 129.360 212.945 130.280 213.175 ;
        RECT 129.360 212.265 132.825 212.945 ;
        RECT 132.945 212.265 134.775 212.945 ;
        RECT 134.785 212.265 138.455 213.075 ;
        RECT 138.465 212.265 139.835 213.075 ;
        RECT 142.500 212.945 143.420 213.175 ;
        RECT 139.955 212.265 143.420 212.945 ;
        RECT 144.455 212.350 144.885 213.135 ;
        RECT 144.905 212.265 146.275 213.045 ;
        RECT 146.285 212.265 147.655 213.045 ;
        RECT 147.665 212.265 151.335 213.075 ;
        RECT 152.265 212.265 153.635 213.045 ;
        RECT 153.645 212.265 156.395 213.075 ;
        RECT 156.865 212.265 158.235 213.075 ;
        RECT 2.905 212.055 3.075 212.265 ;
        RECT 4.285 212.055 4.455 212.265 ;
        RECT 7.965 212.055 8.135 212.245 ;
        RECT 9.805 212.075 9.975 212.265 ;
        RECT 15.320 212.105 15.440 212.215 ;
        RECT 16.245 212.055 16.415 212.265 ;
        RECT 16.700 212.105 16.820 212.215 ;
        RECT 17.165 212.055 17.335 212.245 ;
        RECT 20.845 212.055 21.015 212.245 ;
        RECT 21.765 212.075 21.935 212.265 ;
        RECT 26.365 212.055 26.535 212.245 ;
        RECT 27.285 212.075 27.455 212.265 ;
        RECT 28.200 212.105 28.320 212.215 ;
        RECT 29.125 212.055 29.295 212.245 ;
        RECT 32.805 212.075 32.975 212.265 ;
        RECT 34.645 212.055 34.815 212.245 ;
        RECT 38.325 212.075 38.495 212.265 ;
        RECT 40.165 212.055 40.335 212.245 ;
        RECT 41.080 212.105 41.200 212.215 ;
        RECT 42.005 212.075 42.175 212.265 ;
        RECT 45.685 212.055 45.855 212.245 ;
        RECT 47.525 212.075 47.695 212.265 ;
        RECT 51.205 212.055 51.375 212.245 ;
        RECT 53.045 212.075 53.215 212.265 ;
        RECT 53.960 212.105 54.080 212.215 ;
        RECT 54.885 212.055 55.055 212.245 ;
        RECT 56.725 212.215 56.895 212.265 ;
        RECT 56.720 212.105 56.895 212.215 ;
        RECT 56.725 212.075 56.895 212.105 ;
        RECT 2.765 211.245 4.135 212.055 ;
        RECT 4.145 211.245 7.815 212.055 ;
        RECT 7.825 211.245 9.195 212.055 ;
        RECT 9.245 211.375 16.555 212.055 ;
        RECT 17.135 211.375 20.600 212.055 ;
        RECT 9.245 211.145 10.595 211.375 ;
        RECT 12.130 211.155 13.040 211.375 ;
        RECT 19.680 211.145 20.600 211.375 ;
        RECT 20.705 211.245 26.215 212.055 ;
        RECT 26.225 211.245 28.055 212.055 ;
        RECT 28.535 211.185 28.965 211.970 ;
        RECT 28.985 211.245 34.495 212.055 ;
        RECT 34.505 211.245 40.015 212.055 ;
        RECT 40.025 211.245 45.535 212.055 ;
        RECT 45.545 211.245 51.055 212.055 ;
        RECT 51.065 211.245 53.815 212.055 ;
        RECT 54.295 211.185 54.725 211.970 ;
        RECT 54.745 211.245 56.575 212.055 ;
        RECT 57.190 212.025 57.360 212.245 ;
        RECT 59.485 212.075 59.655 212.265 ;
        RECT 64.085 212.075 64.255 212.265 ;
        RECT 64.545 212.055 64.715 212.265 ;
        RECT 65.010 212.055 65.180 212.245 ;
        RECT 69.145 212.055 69.315 212.245 ;
        RECT 59.320 212.025 60.255 212.055 ;
        RECT 57.190 211.825 60.255 212.025 ;
        RECT 60.275 212.015 61.195 212.055 ;
        RECT 57.045 211.345 60.255 211.825 ;
        RECT 60.265 211.825 61.195 212.015 ;
        RECT 63.285 211.825 64.855 212.055 ;
        RECT 60.265 211.465 64.855 211.825 ;
        RECT 57.045 211.145 57.975 211.345 ;
        RECT 59.305 211.145 60.255 211.345 ;
        RECT 60.275 211.375 64.855 211.465 ;
        RECT 64.865 211.375 68.860 212.055 ;
        RECT 60.275 211.145 63.275 211.375 ;
        RECT 65.350 211.145 68.860 211.375 ;
        RECT 69.005 211.245 70.375 212.055 ;
        RECT 70.530 212.025 70.700 212.245 ;
        RECT 71.440 212.075 71.610 212.265 ;
        RECT 71.905 212.075 72.075 212.265 ;
        RECT 73.750 212.075 73.920 212.265 ;
        RECT 74.205 212.055 74.375 212.245 ;
        RECT 76.050 212.055 76.220 212.245 ;
        RECT 81.560 212.075 81.730 212.265 ;
        RECT 82.485 212.075 82.655 212.245 ;
        RECT 82.485 212.055 82.635 212.075 ;
        RECT 86.620 212.055 86.790 212.245 ;
        RECT 87.085 212.055 87.255 212.245 ;
        RECT 90.765 212.075 90.935 212.265 ;
        RECT 92.605 212.055 92.775 212.265 ;
        RECT 93.525 212.075 93.695 212.265 ;
        RECT 96.295 212.100 96.455 212.210 ;
        RECT 97.205 212.075 97.375 212.245 ;
        RECT 99.045 212.075 99.215 212.265 ;
        RECT 97.225 212.055 97.375 212.075 ;
        RECT 100.425 212.055 100.595 212.245 ;
        RECT 100.885 212.055 101.055 212.245 ;
        RECT 101.800 212.105 101.920 212.215 ;
        RECT 102.540 212.075 102.710 212.265 ;
        RECT 102.725 212.075 102.895 212.245 ;
        RECT 102.745 212.055 102.895 212.075 ;
        RECT 106.405 212.055 106.575 212.245 ;
        RECT 109.625 212.075 109.795 212.265 ;
        RECT 73.105 212.025 74.055 212.055 ;
        RECT 70.385 211.345 74.055 212.025 ;
        RECT 73.105 211.145 74.055 211.345 ;
        RECT 74.065 211.245 75.895 212.055 ;
        RECT 75.905 211.145 79.795 212.055 ;
        RECT 80.055 211.185 80.485 211.970 ;
        RECT 80.705 211.235 82.635 212.055 ;
        RECT 80.705 211.145 81.655 211.235 ;
        RECT 82.900 211.145 86.935 212.055 ;
        RECT 86.945 211.245 92.455 212.055 ;
        RECT 92.465 211.245 96.135 212.055 ;
        RECT 97.225 211.235 99.155 212.055 ;
        RECT 99.365 211.275 100.735 212.055 ;
        RECT 100.745 211.375 102.575 212.055 ;
        RECT 102.745 211.235 104.675 212.055 ;
        RECT 98.205 211.145 99.155 211.235 ;
        RECT 103.725 211.145 104.675 211.235 ;
        RECT 105.815 211.185 106.245 211.970 ;
        RECT 106.275 211.145 109.005 212.055 ;
        RECT 109.025 212.025 110.420 212.055 ;
        RECT 111.465 212.025 111.635 212.245 ;
        RECT 112.840 212.055 113.010 212.245 ;
        RECT 113.305 212.215 113.475 212.265 ;
        RECT 113.300 212.105 113.475 212.215 ;
        RECT 113.305 212.075 113.475 212.105 ;
        RECT 113.765 212.245 113.965 212.265 ;
        RECT 113.765 212.075 113.935 212.245 ;
        RECT 113.765 212.055 113.965 212.075 ;
        RECT 117.445 212.055 117.615 212.245 ;
        RECT 118.365 212.075 118.535 212.265 ;
        RECT 121.125 212.055 121.295 212.245 ;
        RECT 121.585 212.075 121.755 212.265 ;
        RECT 122.045 212.075 122.215 212.265 ;
        RECT 122.505 212.055 122.675 212.245 ;
        RECT 129.865 212.055 130.035 212.245 ;
        RECT 132.625 212.075 132.795 212.265 ;
        RECT 134.465 212.075 134.635 212.265 ;
        RECT 134.925 212.075 135.095 212.265 ;
        RECT 135.385 212.055 135.555 212.245 ;
        RECT 135.845 212.055 136.015 212.245 ;
        RECT 138.605 212.075 138.775 212.265 ;
        RECT 139.985 212.075 140.155 212.265 ;
        RECT 141.365 212.055 141.535 212.245 ;
        RECT 143.675 212.110 143.835 212.220 ;
        RECT 145.045 212.075 145.215 212.265 ;
        RECT 146.885 212.055 147.055 212.245 ;
        RECT 147.345 212.075 147.515 212.265 ;
        RECT 147.805 212.075 147.975 212.265 ;
        RECT 151.495 212.110 151.655 212.220 ;
        RECT 152.405 212.055 152.575 212.245 ;
        RECT 153.325 212.075 153.495 212.265 ;
        RECT 153.785 212.075 153.955 212.265 ;
        RECT 156.095 212.100 156.255 212.210 ;
        RECT 156.540 212.105 156.660 212.215 ;
        RECT 157.925 212.055 158.095 212.265 ;
        RECT 109.025 211.345 111.760 212.025 ;
        RECT 109.025 211.145 110.435 211.345 ;
        RECT 111.805 211.145 113.155 212.055 ;
        RECT 113.765 211.375 117.295 212.055 ;
        RECT 114.470 211.145 117.295 211.375 ;
        RECT 117.305 211.245 120.975 212.055 ;
        RECT 120.985 211.245 122.355 212.055 ;
        RECT 122.365 211.375 129.675 212.055 ;
        RECT 125.880 211.155 126.790 211.375 ;
        RECT 128.325 211.145 129.675 211.375 ;
        RECT 129.725 211.245 131.555 212.055 ;
        RECT 131.575 211.185 132.005 211.970 ;
        RECT 132.120 211.375 135.585 212.055 ;
        RECT 132.120 211.145 133.040 211.375 ;
        RECT 135.705 211.245 141.215 212.055 ;
        RECT 141.225 211.245 146.735 212.055 ;
        RECT 146.745 211.245 152.255 212.055 ;
        RECT 152.265 211.245 155.935 212.055 ;
        RECT 156.865 211.245 158.235 212.055 ;
      LAYER nwell ;
        RECT 2.570 208.025 158.430 210.855 ;
      LAYER pwell ;
        RECT 2.765 206.825 4.135 207.635 ;
        RECT 4.145 206.825 9.655 207.635 ;
        RECT 14.620 207.505 15.540 207.735 ;
        RECT 12.075 206.825 15.540 207.505 ;
        RECT 15.655 206.910 16.085 207.695 ;
        RECT 16.105 206.825 18.855 207.635 ;
        RECT 22.840 207.505 23.750 207.725 ;
        RECT 25.285 207.505 27.055 207.735 ;
        RECT 19.325 206.825 27.055 207.505 ;
        RECT 27.145 206.825 29.895 207.635 ;
        RECT 32.560 207.505 33.480 207.735 ;
        RECT 30.015 206.825 33.480 207.505 ;
        RECT 33.585 206.825 39.095 207.635 ;
        RECT 39.105 206.825 40.935 207.635 ;
        RECT 41.415 206.910 41.845 207.695 ;
        RECT 41.865 206.825 47.375 207.635 ;
        RECT 47.385 206.825 52.895 207.635 ;
        RECT 52.905 206.825 58.415 207.635 ;
        RECT 58.665 206.825 62.555 207.735 ;
        RECT 62.805 206.825 66.695 207.735 ;
        RECT 67.175 206.910 67.605 207.695 ;
        RECT 67.635 206.825 68.985 207.735 ;
        RECT 69.465 206.825 76.815 207.735 ;
        RECT 77.965 207.645 78.915 207.735 ;
        RECT 76.985 206.825 78.915 207.645 ;
        RECT 79.125 206.825 80.495 207.635 ;
        RECT 80.640 207.505 84.150 207.735 ;
        RECT 85.785 207.645 86.735 207.735 ;
        RECT 90.845 207.645 91.795 207.735 ;
        RECT 80.640 206.825 84.635 207.505 ;
        RECT 84.805 206.825 86.735 207.645 ;
        RECT 86.945 206.825 89.695 207.635 ;
        RECT 89.865 206.825 91.795 207.645 ;
        RECT 92.935 206.910 93.365 207.695 ;
        RECT 97.285 207.645 98.235 207.735 ;
        RECT 93.385 206.825 96.135 207.635 ;
        RECT 96.305 206.825 98.235 207.645 ;
        RECT 102.955 207.505 103.885 207.725 ;
        RECT 106.605 207.505 108.815 207.735 ;
        RECT 98.445 206.825 108.815 207.505 ;
        RECT 109.225 207.645 110.175 207.735 ;
        RECT 109.225 206.825 111.155 207.645 ;
        RECT 111.405 206.825 113.615 207.735 ;
        RECT 113.625 206.825 117.295 207.635 ;
        RECT 117.305 206.825 118.675 207.635 ;
        RECT 118.695 206.910 119.125 207.695 ;
        RECT 119.145 206.825 124.655 207.635 ;
        RECT 124.665 206.825 126.495 207.635 ;
        RECT 128.770 207.535 129.715 207.735 ;
        RECT 126.965 206.855 129.715 207.535 ;
        RECT 2.905 206.615 3.075 206.825 ;
        RECT 4.285 206.615 4.455 206.825 ;
        RECT 9.815 206.775 9.975 206.780 ;
        RECT 9.800 206.670 9.975 206.775 ;
        RECT 9.800 206.665 9.920 206.670 ;
        RECT 11.645 206.615 11.815 206.805 ;
        RECT 12.105 206.635 12.275 206.825 ;
        RECT 16.245 206.635 16.415 206.825 ;
        RECT 19.000 206.665 19.120 206.775 ;
        RECT 19.465 206.615 19.635 206.825 ;
        RECT 19.925 206.615 20.095 206.805 ;
        RECT 22.685 206.615 22.855 206.805 ;
        RECT 23.145 206.615 23.315 206.805 ;
        RECT 27.285 206.635 27.455 206.825 ;
        RECT 29.125 206.615 29.295 206.805 ;
        RECT 30.045 206.635 30.215 206.825 ;
        RECT 31.880 206.665 32.000 206.775 ;
        RECT 33.725 206.615 33.895 206.825 ;
        RECT 34.185 206.615 34.355 206.805 ;
        RECT 39.245 206.635 39.415 206.825 ;
        RECT 41.085 206.775 41.255 206.805 ;
        RECT 41.080 206.665 41.255 206.775 ;
        RECT 41.085 206.615 41.255 206.665 ;
        RECT 41.545 206.615 41.715 206.805 ;
        RECT 42.005 206.635 42.175 206.825 ;
        RECT 47.065 206.615 47.235 206.805 ;
        RECT 47.525 206.635 47.695 206.825 ;
        RECT 52.585 206.615 52.755 206.805 ;
        RECT 53.045 206.635 53.215 206.825 ;
        RECT 54.885 206.615 55.055 206.805 ;
        RECT 58.570 206.615 58.740 206.805 ;
        RECT 62.240 206.635 62.410 206.825 ;
        RECT 66.380 206.635 66.550 206.825 ;
        RECT 66.840 206.665 66.960 206.775 ;
        RECT 68.220 206.615 68.390 206.805 ;
        RECT 68.685 206.635 68.855 206.825 ;
        RECT 69.140 206.665 69.260 206.775 ;
        RECT 71.440 206.615 71.610 206.805 ;
        RECT 75.580 206.615 75.750 206.805 ;
        RECT 76.500 206.635 76.670 206.825 ;
        RECT 76.985 206.805 77.135 206.825 ;
        RECT 76.965 206.635 77.135 206.805 ;
        RECT 79.265 206.635 79.435 206.825 ;
        RECT 79.720 206.615 79.890 206.805 ;
        RECT 84.320 206.615 84.490 206.825 ;
        RECT 84.805 206.805 84.955 206.825 ;
        RECT 84.785 206.635 84.960 206.805 ;
        RECT 87.085 206.635 87.255 206.825 ;
        RECT 89.865 206.805 90.015 206.825 ;
        RECT 84.790 206.615 84.960 206.635 ;
        RECT 88.925 206.615 89.095 206.805 ;
        RECT 89.845 206.635 90.015 206.805 ;
        RECT 90.765 206.615 90.935 206.805 ;
        RECT 92.155 206.670 92.315 206.780 ;
        RECT 93.525 206.635 93.695 206.825 ;
        RECT 96.305 206.805 96.455 206.825 ;
        RECT 94.445 206.615 94.615 206.805 ;
        RECT 95.825 206.615 95.995 206.805 ;
        RECT 96.285 206.635 96.455 206.805 ;
        RECT 98.585 206.615 98.755 206.825 ;
        RECT 111.005 206.805 111.155 206.825 ;
        RECT 101.345 206.615 101.515 206.805 ;
        RECT 103.185 206.615 103.355 206.805 ;
        RECT 106.415 206.660 106.575 206.770 ;
        RECT 109.625 206.615 109.795 206.805 ;
        RECT 110.085 206.615 110.255 206.805 ;
        RECT 111.005 206.635 111.175 206.805 ;
        RECT 111.925 206.615 112.095 206.805 ;
        RECT 113.300 206.635 113.470 206.825 ;
        RECT 113.765 206.635 113.935 206.825 ;
        RECT 117.445 206.615 117.615 206.825 ;
        RECT 118.825 206.615 118.995 206.805 ;
        RECT 119.285 206.635 119.455 206.825 ;
        RECT 124.345 206.615 124.515 206.805 ;
        RECT 124.805 206.635 124.975 206.825 ;
        RECT 126.640 206.665 126.760 206.775 ;
        RECT 127.110 206.635 127.280 206.855 ;
        RECT 128.770 206.825 129.715 206.855 ;
        RECT 129.725 206.825 135.235 207.635 ;
        RECT 135.245 206.825 140.755 207.635 ;
        RECT 140.765 206.825 144.435 207.635 ;
        RECT 144.455 206.910 144.885 207.695 ;
        RECT 144.905 206.825 150.415 207.635 ;
        RECT 150.425 206.825 155.935 207.635 ;
        RECT 156.865 206.825 158.235 207.635 ;
        RECT 129.865 206.615 130.035 206.825 ;
        RECT 132.165 206.615 132.335 206.805 ;
        RECT 135.385 206.635 135.555 206.825 ;
        RECT 137.685 206.615 137.855 206.805 ;
        RECT 140.905 206.635 141.075 206.825 ;
        RECT 143.205 206.615 143.375 206.805 ;
        RECT 145.045 206.635 145.215 206.825 ;
        RECT 148.725 206.615 148.895 206.805 ;
        RECT 150.565 206.635 150.735 206.825 ;
        RECT 152.400 206.615 152.570 206.805 ;
        RECT 152.865 206.615 153.035 206.805 ;
        RECT 156.095 206.670 156.255 206.780 ;
        RECT 156.540 206.665 156.660 206.775 ;
        RECT 157.925 206.615 158.095 206.825 ;
        RECT 2.765 205.805 4.135 206.615 ;
        RECT 4.145 205.805 9.655 206.615 ;
        RECT 10.125 205.935 11.955 206.615 ;
        RECT 12.045 205.935 19.775 206.615 ;
        RECT 10.125 205.705 11.470 205.935 ;
        RECT 12.045 205.705 13.815 205.935 ;
        RECT 15.350 205.715 16.260 205.935 ;
        RECT 19.785 205.805 21.155 206.615 ;
        RECT 21.165 205.935 22.995 206.615 ;
        RECT 21.165 205.705 22.510 205.935 ;
        RECT 23.005 205.805 28.515 206.615 ;
        RECT 28.535 205.745 28.965 206.530 ;
        RECT 28.985 205.805 31.735 206.615 ;
        RECT 32.205 205.935 34.035 206.615 ;
        RECT 32.205 205.705 33.550 205.935 ;
        RECT 34.045 205.805 39.555 206.615 ;
        RECT 39.565 205.935 41.395 206.615 ;
        RECT 39.565 205.705 40.910 205.935 ;
        RECT 41.405 205.805 46.915 206.615 ;
        RECT 46.925 205.805 52.435 206.615 ;
        RECT 52.445 205.805 54.275 206.615 ;
        RECT 54.295 205.745 54.725 206.530 ;
        RECT 54.745 205.805 58.415 206.615 ;
        RECT 58.425 205.705 62.315 206.615 ;
        RECT 62.965 205.705 68.535 206.615 ;
        RECT 68.640 205.705 71.755 206.615 ;
        RECT 72.005 205.705 75.895 206.615 ;
        RECT 76.145 205.705 80.035 206.615 ;
        RECT 80.055 205.745 80.485 206.530 ;
        RECT 80.745 205.705 84.635 206.615 ;
        RECT 84.645 205.705 88.535 206.615 ;
        RECT 88.785 205.935 90.615 206.615 ;
        RECT 89.270 205.705 90.615 205.935 ;
        RECT 90.625 205.805 94.295 206.615 ;
        RECT 94.305 205.805 95.675 206.615 ;
        RECT 95.685 205.935 98.425 206.615 ;
        RECT 98.445 205.805 101.195 206.615 ;
        RECT 101.205 205.935 103.035 206.615 ;
        RECT 103.045 205.935 105.785 206.615 ;
        RECT 101.690 205.705 103.035 205.935 ;
        RECT 105.815 205.745 106.245 206.530 ;
        RECT 107.195 205.935 109.935 206.615 ;
        RECT 109.945 205.935 111.775 206.615 ;
        RECT 110.430 205.705 111.775 205.935 ;
        RECT 111.785 205.805 117.295 206.615 ;
        RECT 117.315 205.705 118.665 206.615 ;
        RECT 118.685 205.805 124.195 206.615 ;
        RECT 124.205 205.805 129.715 206.615 ;
        RECT 129.725 205.805 131.555 206.615 ;
        RECT 131.575 205.745 132.005 206.530 ;
        RECT 132.025 205.805 137.535 206.615 ;
        RECT 137.545 205.805 143.055 206.615 ;
        RECT 143.065 205.805 148.575 206.615 ;
        RECT 148.585 205.805 149.955 206.615 ;
        RECT 150.105 205.705 152.715 206.615 ;
        RECT 152.725 205.805 156.395 206.615 ;
        RECT 156.865 205.805 158.235 206.615 ;
      LAYER nwell ;
        RECT 2.570 202.585 158.430 205.415 ;
      LAYER pwell ;
        RECT 2.765 201.385 4.135 202.195 ;
        RECT 4.145 201.385 9.655 202.195 ;
        RECT 9.665 201.385 15.175 202.195 ;
        RECT 15.655 201.470 16.085 202.255 ;
        RECT 16.105 201.385 21.615 202.195 ;
        RECT 21.625 201.385 27.135 202.195 ;
        RECT 27.145 201.385 28.515 202.195 ;
        RECT 28.535 201.470 28.965 202.255 ;
        RECT 28.985 201.385 34.495 202.195 ;
        RECT 34.505 201.385 40.015 202.195 ;
        RECT 40.025 201.385 41.395 202.195 ;
        RECT 41.415 201.470 41.845 202.255 ;
        RECT 41.865 201.385 47.375 202.195 ;
        RECT 47.385 201.385 52.895 202.195 ;
        RECT 52.905 201.385 54.275 202.195 ;
        RECT 54.295 201.470 54.725 202.255 ;
        RECT 63.685 202.205 64.635 202.295 ;
        RECT 54.745 201.385 60.255 202.195 ;
        RECT 60.265 201.385 63.015 202.195 ;
        RECT 63.685 201.385 65.615 202.205 ;
        RECT 65.785 201.385 67.155 202.195 ;
        RECT 67.175 201.470 67.605 202.255 ;
        RECT 67.625 201.385 73.135 202.195 ;
        RECT 73.145 201.385 74.975 202.195 ;
        RECT 75.225 201.385 79.115 202.295 ;
        RECT 80.055 201.470 80.485 202.255 ;
        RECT 80.990 202.065 82.335 202.295 ;
        RECT 80.505 201.385 82.335 202.065 ;
        RECT 82.345 201.385 87.855 202.195 ;
        RECT 87.865 201.385 91.535 202.195 ;
        RECT 91.545 201.385 92.915 202.195 ;
        RECT 92.935 201.470 93.365 202.255 ;
        RECT 93.385 201.385 98.895 202.195 ;
        RECT 98.905 201.385 104.415 202.195 ;
        RECT 104.425 201.385 105.795 202.195 ;
        RECT 105.815 201.470 106.245 202.255 ;
        RECT 106.265 201.385 111.775 202.195 ;
        RECT 111.785 201.385 117.295 202.195 ;
        RECT 117.305 201.385 118.675 202.195 ;
        RECT 118.695 201.470 119.125 202.255 ;
        RECT 119.145 201.385 124.655 202.195 ;
        RECT 124.665 201.385 130.175 202.195 ;
        RECT 130.185 201.385 131.555 202.195 ;
        RECT 131.575 201.470 132.005 202.255 ;
        RECT 132.025 201.385 137.535 202.195 ;
        RECT 137.545 201.385 143.055 202.195 ;
        RECT 143.065 201.385 144.435 202.195 ;
        RECT 144.455 201.470 144.885 202.255 ;
        RECT 144.905 201.385 150.415 202.195 ;
        RECT 150.425 201.385 155.935 202.195 ;
        RECT 156.865 201.385 158.235 202.195 ;
        RECT 2.905 201.195 3.075 201.385 ;
        RECT 4.285 201.195 4.455 201.385 ;
        RECT 9.805 201.195 9.975 201.385 ;
        RECT 15.320 201.225 15.440 201.335 ;
        RECT 16.245 201.195 16.415 201.385 ;
        RECT 21.765 201.195 21.935 201.385 ;
        RECT 27.285 201.195 27.455 201.385 ;
        RECT 29.125 201.195 29.295 201.385 ;
        RECT 34.645 201.195 34.815 201.385 ;
        RECT 40.165 201.195 40.335 201.385 ;
        RECT 42.005 201.195 42.175 201.385 ;
        RECT 47.525 201.195 47.695 201.385 ;
        RECT 53.045 201.195 53.215 201.385 ;
        RECT 54.885 201.195 55.055 201.385 ;
        RECT 60.405 201.195 60.575 201.385 ;
        RECT 65.465 201.365 65.615 201.385 ;
        RECT 63.160 201.225 63.280 201.335 ;
        RECT 65.465 201.195 65.635 201.365 ;
        RECT 65.925 201.195 66.095 201.385 ;
        RECT 67.765 201.195 67.935 201.385 ;
        RECT 73.285 201.195 73.455 201.385 ;
        RECT 78.800 201.195 78.970 201.385 ;
        RECT 79.275 201.230 79.435 201.340 ;
        RECT 80.645 201.195 80.815 201.385 ;
        RECT 82.485 201.195 82.655 201.385 ;
        RECT 88.005 201.195 88.175 201.385 ;
        RECT 91.685 201.195 91.855 201.385 ;
        RECT 93.525 201.195 93.695 201.385 ;
        RECT 99.045 201.195 99.215 201.385 ;
        RECT 104.565 201.195 104.735 201.385 ;
        RECT 106.405 201.195 106.575 201.385 ;
        RECT 111.925 201.195 112.095 201.385 ;
        RECT 117.445 201.195 117.615 201.385 ;
        RECT 119.285 201.195 119.455 201.385 ;
        RECT 124.805 201.195 124.975 201.385 ;
        RECT 130.325 201.195 130.495 201.385 ;
        RECT 132.165 201.195 132.335 201.385 ;
        RECT 137.685 201.195 137.855 201.385 ;
        RECT 143.205 201.195 143.375 201.385 ;
        RECT 145.045 201.195 145.215 201.385 ;
        RECT 150.565 201.195 150.735 201.385 ;
        RECT 156.095 201.230 156.255 201.340 ;
        RECT 157.925 201.195 158.095 201.385 ;
        RECT 2.800 197.810 93.920 199.820 ;
      LAYER nwell ;
        RECT 10.600 158.310 19.310 166.500 ;
        RECT 17.200 156.500 19.310 158.310 ;
        RECT 10.600 148.310 19.310 156.500 ;
      LAYER pwell ;
        RECT 20.560 158.310 25.430 164.410 ;
        RECT 20.560 156.020 22.670 158.310 ;
        RECT 23.200 156.010 25.310 158.310 ;
      LAYER nwell ;
        RECT 134.140 158.300 142.850 166.490 ;
        RECT 140.740 156.490 142.850 158.300 ;
        RECT 17.200 146.500 19.310 148.310 ;
        RECT 10.600 138.310 19.310 146.500 ;
      LAYER pwell ;
        RECT 20.560 148.310 25.430 154.410 ;
        RECT 20.560 146.020 22.670 148.310 ;
        RECT 23.200 146.010 25.310 148.310 ;
      LAYER nwell ;
        RECT 134.140 148.300 142.850 156.490 ;
      LAYER pwell ;
        RECT 144.100 158.300 148.970 164.400 ;
        RECT 144.100 156.010 146.210 158.300 ;
      LAYER nwell ;
        RECT 140.740 146.490 142.850 148.300 ;
        RECT 17.200 136.500 19.310 138.310 ;
        RECT 10.600 128.310 19.310 136.500 ;
      LAYER pwell ;
        RECT 20.560 138.310 25.430 144.410 ;
        RECT 20.560 136.020 22.670 138.310 ;
        RECT 23.200 136.010 25.310 138.310 ;
      LAYER nwell ;
        RECT 134.140 138.300 142.850 146.490 ;
      LAYER pwell ;
        RECT 144.100 148.300 148.970 154.400 ;
        RECT 144.100 146.010 146.210 148.300 ;
      LAYER nwell ;
        RECT 140.740 136.490 142.850 138.300 ;
        RECT 17.200 126.500 19.310 128.310 ;
        RECT 10.600 118.310 19.310 126.500 ;
      LAYER pwell ;
        RECT 20.560 128.310 25.430 134.410 ;
        RECT 20.560 126.020 22.670 128.310 ;
        RECT 23.200 126.010 25.310 128.310 ;
      LAYER nwell ;
        RECT 134.140 128.300 142.850 136.490 ;
      LAYER pwell ;
        RECT 144.100 138.300 148.970 144.400 ;
        RECT 144.100 136.010 146.210 138.300 ;
      LAYER nwell ;
        RECT 140.740 126.490 142.850 128.300 ;
        RECT 17.200 116.500 19.310 118.310 ;
        RECT 10.600 108.310 19.310 116.500 ;
      LAYER pwell ;
        RECT 20.560 118.310 25.430 124.410 ;
        RECT 20.560 116.020 22.670 118.310 ;
        RECT 23.200 116.010 25.310 118.310 ;
      LAYER nwell ;
        RECT 134.140 118.300 142.850 126.490 ;
      LAYER pwell ;
        RECT 144.100 128.300 148.970 134.400 ;
        RECT 144.100 126.010 146.210 128.300 ;
      LAYER nwell ;
        RECT 140.740 116.490 142.850 118.300 ;
        RECT 17.200 106.500 19.310 108.310 ;
        RECT 10.600 98.310 19.310 106.500 ;
      LAYER pwell ;
        RECT 20.560 108.310 25.430 114.410 ;
        RECT 20.560 106.020 22.670 108.310 ;
        RECT 23.200 106.010 25.310 108.310 ;
      LAYER nwell ;
        RECT 134.140 108.300 142.850 116.490 ;
      LAYER pwell ;
        RECT 144.100 118.300 148.970 124.400 ;
        RECT 144.100 116.010 146.210 118.300 ;
      LAYER nwell ;
        RECT 140.740 106.490 142.850 108.300 ;
        RECT 17.200 96.500 19.310 98.310 ;
        RECT 10.600 88.310 19.310 96.500 ;
      LAYER pwell ;
        RECT 20.560 98.310 25.430 104.410 ;
        RECT 20.560 96.020 22.670 98.310 ;
        RECT 23.200 96.010 25.310 98.310 ;
      LAYER nwell ;
        RECT 134.140 98.300 142.850 106.490 ;
      LAYER pwell ;
        RECT 144.100 108.300 148.970 114.400 ;
        RECT 144.100 106.010 146.210 108.300 ;
      LAYER nwell ;
        RECT 140.740 96.490 142.850 98.300 ;
        RECT 17.200 86.500 19.310 88.310 ;
        RECT 10.600 78.310 19.310 86.500 ;
      LAYER pwell ;
        RECT 20.560 88.310 25.430 94.410 ;
        RECT 20.560 86.020 22.670 88.310 ;
        RECT 23.200 86.010 25.310 88.310 ;
      LAYER nwell ;
        RECT 134.140 88.300 142.850 96.490 ;
      LAYER pwell ;
        RECT 144.100 98.300 148.970 104.400 ;
        RECT 144.100 96.010 146.210 98.300 ;
      LAYER nwell ;
        RECT 140.740 86.490 142.850 88.300 ;
        RECT 17.200 76.500 19.310 78.310 ;
        RECT 10.600 68.310 19.310 76.500 ;
      LAYER pwell ;
        RECT 20.560 78.310 25.430 84.410 ;
        RECT 20.560 76.020 22.670 78.310 ;
        RECT 23.200 76.010 25.310 78.310 ;
      LAYER nwell ;
        RECT 134.140 78.300 142.850 86.490 ;
      LAYER pwell ;
        RECT 144.100 88.300 148.970 94.400 ;
        RECT 144.100 86.010 146.210 88.300 ;
      LAYER nwell ;
        RECT 140.740 76.490 142.850 78.300 ;
        RECT 17.200 66.500 19.310 68.310 ;
        RECT 10.600 58.310 19.310 66.500 ;
      LAYER pwell ;
        RECT 20.560 68.310 25.430 74.410 ;
        RECT 20.560 66.020 22.670 68.310 ;
        RECT 23.200 66.010 25.310 68.310 ;
      LAYER nwell ;
        RECT 134.140 68.300 142.850 76.490 ;
      LAYER pwell ;
        RECT 144.100 78.300 148.970 84.400 ;
        RECT 144.100 76.010 146.210 78.300 ;
      LAYER nwell ;
        RECT 140.740 66.490 142.850 68.300 ;
        RECT 17.200 56.500 19.310 58.310 ;
        RECT 10.600 48.310 19.310 56.500 ;
      LAYER pwell ;
        RECT 20.560 58.310 25.430 64.410 ;
        RECT 20.560 56.020 22.670 58.310 ;
        RECT 23.200 56.010 25.310 58.310 ;
      LAYER nwell ;
        RECT 134.140 58.300 142.850 66.490 ;
      LAYER pwell ;
        RECT 144.100 68.300 148.970 74.400 ;
        RECT 144.100 66.010 146.210 68.300 ;
      LAYER nwell ;
        RECT 140.740 56.490 142.850 58.300 ;
        RECT 17.200 46.500 19.310 48.310 ;
        RECT 10.600 38.310 19.310 46.500 ;
      LAYER pwell ;
        RECT 20.560 48.310 25.430 54.410 ;
        RECT 20.560 46.020 22.670 48.310 ;
        RECT 23.200 46.010 25.310 48.310 ;
      LAYER nwell ;
        RECT 134.140 48.300 142.850 56.490 ;
      LAYER pwell ;
        RECT 144.100 58.300 148.970 64.400 ;
        RECT 144.100 56.010 146.210 58.300 ;
      LAYER nwell ;
        RECT 140.740 46.490 142.850 48.300 ;
        RECT 17.200 36.500 19.310 38.310 ;
        RECT 10.600 28.310 19.310 36.500 ;
      LAYER pwell ;
        RECT 20.560 38.310 25.430 44.410 ;
        RECT 20.560 36.020 22.670 38.310 ;
        RECT 23.200 36.010 25.310 38.310 ;
      LAYER nwell ;
        RECT 134.140 38.300 142.850 46.490 ;
      LAYER pwell ;
        RECT 144.100 48.300 148.970 54.400 ;
        RECT 144.100 46.010 146.210 48.300 ;
      LAYER nwell ;
        RECT 140.740 36.490 142.850 38.300 ;
        RECT 17.200 26.500 19.310 28.310 ;
        RECT 10.600 18.310 19.310 26.500 ;
      LAYER pwell ;
        RECT 20.560 28.310 25.430 34.410 ;
        RECT 20.560 26.020 22.670 28.310 ;
        RECT 23.200 26.010 25.310 28.310 ;
      LAYER nwell ;
        RECT 134.140 28.300 142.850 36.490 ;
      LAYER pwell ;
        RECT 144.100 38.300 148.970 44.400 ;
        RECT 144.100 36.010 146.210 38.300 ;
      LAYER nwell ;
        RECT 140.740 26.490 142.850 28.300 ;
        RECT 17.200 16.500 19.310 18.310 ;
        RECT 10.600 8.310 19.310 16.500 ;
      LAYER pwell ;
        RECT 20.560 18.310 25.430 24.410 ;
        RECT 20.560 16.020 22.670 18.310 ;
        RECT 23.200 16.010 25.310 18.310 ;
      LAYER nwell ;
        RECT 134.140 18.300 142.850 26.490 ;
      LAYER pwell ;
        RECT 144.100 28.300 148.970 34.400 ;
        RECT 144.100 26.010 146.210 28.300 ;
      LAYER nwell ;
        RECT 140.740 16.490 142.850 18.300 ;
        RECT 17.200 6.000 19.310 8.310 ;
      LAYER pwell ;
        RECT 20.560 8.310 25.430 14.410 ;
        RECT 20.560 6.020 22.670 8.310 ;
        RECT 23.200 6.010 25.310 8.310 ;
      LAYER nwell ;
        RECT 134.140 8.300 142.850 16.490 ;
      LAYER pwell ;
        RECT 144.100 18.300 148.970 24.400 ;
        RECT 144.100 16.010 146.210 18.300 ;
      LAYER nwell ;
        RECT 140.740 5.990 142.850 8.300 ;
      LAYER pwell ;
        RECT 144.100 8.300 148.970 14.400 ;
        RECT 144.100 6.010 146.210 8.300 ;
      LAYER li1 ;
        RECT 2.760 222.955 158.240 223.125 ;
        RECT 2.845 222.205 4.055 222.955 ;
        RECT 2.845 221.665 3.365 222.205 ;
        RECT 3.535 221.495 4.055 222.035 ;
        RECT 2.845 220.405 4.055 221.495 ;
        RECT 4.225 221.300 4.745 222.785 ;
        RECT 4.915 222.295 5.255 222.955 ;
        RECT 5.605 222.185 7.275 222.955 ;
        RECT 4.415 220.405 4.745 221.130 ;
        RECT 4.915 220.575 5.435 222.125 ;
        RECT 5.605 221.665 6.355 222.185 ;
        RECT 6.525 221.495 7.275 222.015 ;
        RECT 5.605 220.405 7.275 221.495 ;
        RECT 7.905 221.300 8.425 222.785 ;
        RECT 8.595 222.295 8.935 222.955 ;
        RECT 9.285 222.185 10.955 222.955 ;
        RECT 8.095 220.405 8.425 221.130 ;
        RECT 8.595 220.575 9.115 222.125 ;
        RECT 9.285 221.665 10.035 222.185 ;
        RECT 10.205 221.495 10.955 222.015 ;
        RECT 9.285 220.405 10.955 221.495 ;
        RECT 11.585 221.300 12.105 222.785 ;
        RECT 12.275 222.295 12.615 222.955 ;
        RECT 12.965 222.185 15.555 222.955 ;
        RECT 15.725 222.230 16.015 222.955 ;
        RECT 11.775 220.405 12.105 221.130 ;
        RECT 12.275 220.575 12.795 222.125 ;
        RECT 12.965 221.665 14.175 222.185 ;
        RECT 14.345 221.495 15.555 222.015 ;
        RECT 12.965 220.405 15.555 221.495 ;
        RECT 15.725 220.405 16.015 221.570 ;
        RECT 16.185 221.300 16.705 222.785 ;
        RECT 16.875 222.295 17.215 222.955 ;
        RECT 17.565 222.205 18.775 222.955 ;
        RECT 16.375 220.405 16.705 221.130 ;
        RECT 16.875 220.575 17.395 222.125 ;
        RECT 17.565 221.665 18.085 222.205 ;
        RECT 18.255 221.495 18.775 222.035 ;
        RECT 17.565 220.405 18.775 221.495 ;
        RECT 18.945 221.300 19.465 222.785 ;
        RECT 19.635 222.295 19.975 222.955 ;
        RECT 20.325 222.185 21.995 222.955 ;
        RECT 19.135 220.405 19.465 221.130 ;
        RECT 19.635 220.575 20.155 222.125 ;
        RECT 20.325 221.665 21.075 222.185 ;
        RECT 21.245 221.495 21.995 222.015 ;
        RECT 20.325 220.405 21.995 221.495 ;
        RECT 22.625 221.300 23.145 222.785 ;
        RECT 23.315 222.295 23.655 222.955 ;
        RECT 24.005 222.185 25.675 222.955 ;
        RECT 22.815 220.405 23.145 221.130 ;
        RECT 23.315 220.575 23.835 222.125 ;
        RECT 24.005 221.665 24.755 222.185 ;
        RECT 24.925 221.495 25.675 222.015 ;
        RECT 24.005 220.405 25.675 221.495 ;
        RECT 26.305 221.300 26.825 222.785 ;
        RECT 26.995 222.295 27.335 222.955 ;
        RECT 28.605 222.230 28.895 222.955 ;
        RECT 26.495 220.405 26.825 221.130 ;
        RECT 26.995 220.575 27.515 222.125 ;
        RECT 28.605 220.405 28.895 221.570 ;
        RECT 29.985 221.300 30.505 222.785 ;
        RECT 30.675 222.295 31.015 222.955 ;
        RECT 31.365 222.410 36.710 222.955 ;
        RECT 30.175 220.405 30.505 221.130 ;
        RECT 30.675 220.575 31.195 222.125 ;
        RECT 32.950 221.580 33.290 222.410 ;
        RECT 36.885 222.185 40.395 222.955 ;
        RECT 41.485 222.230 41.775 222.955 ;
        RECT 41.945 222.410 47.290 222.955 ;
        RECT 47.465 222.410 52.810 222.955 ;
        RECT 34.770 220.840 35.120 222.090 ;
        RECT 36.885 221.665 38.535 222.185 ;
        RECT 38.705 221.495 40.395 222.015 ;
        RECT 43.530 221.580 43.870 222.410 ;
        RECT 31.365 220.405 36.710 220.840 ;
        RECT 36.885 220.405 40.395 221.495 ;
        RECT 41.485 220.405 41.775 221.570 ;
        RECT 45.350 220.840 45.700 222.090 ;
        RECT 49.050 221.580 49.390 222.410 ;
        RECT 52.985 222.205 54.195 222.955 ;
        RECT 54.365 222.230 54.655 222.955 ;
        RECT 50.870 220.840 51.220 222.090 ;
        RECT 52.985 221.665 53.505 222.205 ;
        RECT 54.825 222.185 57.415 222.955 ;
        RECT 58.260 222.485 58.545 222.955 ;
        RECT 58.715 222.315 59.045 222.785 ;
        RECT 59.215 222.485 59.385 222.955 ;
        RECT 59.555 222.315 59.885 222.785 ;
        RECT 60.055 222.485 60.225 222.955 ;
        RECT 60.395 222.315 60.725 222.785 ;
        RECT 60.895 222.485 61.065 222.955 ;
        RECT 61.235 222.315 61.565 222.785 ;
        RECT 53.675 221.495 54.195 222.035 ;
        RECT 54.825 221.665 56.035 222.185 ;
        RECT 58.045 222.135 61.565 222.315 ;
        RECT 61.735 222.135 62.010 222.955 ;
        RECT 62.650 222.700 62.985 222.745 ;
        RECT 62.645 222.235 62.985 222.700 ;
        RECT 63.155 222.575 63.485 222.955 ;
        RECT 41.945 220.405 47.290 220.840 ;
        RECT 47.465 220.405 52.810 220.840 ;
        RECT 52.985 220.405 54.195 221.495 ;
        RECT 54.365 220.405 54.655 221.570 ;
        RECT 56.205 221.495 57.415 222.015 ;
        RECT 54.825 220.405 57.415 221.495 ;
        RECT 58.045 221.595 58.445 222.135 ;
        RECT 58.615 221.765 59.980 221.965 ;
        RECT 60.300 221.765 61.960 221.965 ;
        RECT 58.045 221.295 59.805 221.595 ;
        RECT 58.210 220.745 58.625 221.125 ;
        RECT 58.795 220.915 58.965 221.295 ;
        RECT 59.135 220.745 59.465 221.105 ;
        RECT 59.635 220.915 59.805 221.295 ;
        RECT 59.975 221.375 62.010 221.585 ;
        RECT 59.975 220.745 60.305 221.375 ;
        RECT 58.210 220.575 60.305 220.745 ;
        RECT 60.475 220.405 60.725 221.205 ;
        RECT 60.895 220.575 61.065 221.375 ;
        RECT 61.235 220.405 61.565 221.205 ;
        RECT 61.735 220.575 62.010 221.375 ;
        RECT 62.645 221.545 62.815 222.235 ;
        RECT 62.985 221.715 63.245 222.045 ;
        RECT 62.645 220.575 62.905 221.545 ;
        RECT 63.075 221.165 63.245 221.715 ;
        RECT 63.415 221.345 63.755 222.375 ;
        RECT 63.945 221.505 64.215 222.620 ;
        RECT 63.945 221.345 64.255 221.505 ;
        RECT 64.440 221.345 64.720 222.620 ;
        RECT 64.920 222.455 65.150 222.785 ;
        RECT 65.395 222.575 65.725 222.955 ;
        RECT 63.500 221.335 63.670 221.345 ;
        RECT 64.085 221.335 64.255 221.345 ;
        RECT 64.920 221.165 65.090 222.455 ;
        RECT 65.895 222.385 66.070 222.785 ;
        RECT 65.440 222.215 66.070 222.385 ;
        RECT 67.245 222.230 67.535 222.955 ;
        RECT 67.815 222.575 68.985 222.785 ;
        RECT 67.815 222.555 68.145 222.575 ;
        RECT 65.440 222.045 65.610 222.215 ;
        RECT 67.705 222.135 68.565 222.385 ;
        RECT 68.735 222.325 68.985 222.575 ;
        RECT 69.155 222.495 69.325 222.955 ;
        RECT 69.495 222.325 69.835 222.785 ;
        RECT 68.735 222.155 69.835 222.325 ;
        RECT 65.260 221.715 65.610 222.045 ;
        RECT 63.075 220.995 65.090 221.165 ;
        RECT 65.440 221.195 65.610 221.715 ;
        RECT 65.790 221.365 66.155 222.045 ;
        RECT 65.440 221.025 66.070 221.195 ;
        RECT 63.100 220.405 63.430 220.815 ;
        RECT 63.630 220.575 63.800 220.995 ;
        RECT 64.015 220.405 64.685 220.815 ;
        RECT 64.920 220.575 65.090 220.995 ;
        RECT 65.395 220.405 65.725 220.845 ;
        RECT 65.895 220.575 66.070 221.025 ;
        RECT 67.245 220.405 67.535 221.570 ;
        RECT 67.705 221.545 67.985 222.135 ;
        RECT 70.010 222.115 70.270 222.955 ;
        RECT 70.445 222.210 70.700 222.785 ;
        RECT 70.870 222.575 71.200 222.955 ;
        RECT 71.415 222.405 71.585 222.785 ;
        RECT 71.845 222.410 77.190 222.955 ;
        RECT 70.870 222.235 71.585 222.405 ;
        RECT 68.155 221.715 68.905 221.965 ;
        RECT 69.075 221.715 69.835 221.965 ;
        RECT 67.705 221.375 69.405 221.545 ;
        RECT 67.810 220.405 68.065 221.205 ;
        RECT 68.235 220.575 68.565 221.375 ;
        RECT 68.735 220.405 68.905 221.205 ;
        RECT 69.075 220.575 69.405 221.375 ;
        RECT 69.575 220.405 69.835 221.545 ;
        RECT 70.010 220.405 70.270 221.555 ;
        RECT 70.445 221.480 70.615 222.210 ;
        RECT 70.870 222.045 71.040 222.235 ;
        RECT 70.785 221.715 71.040 222.045 ;
        RECT 70.870 221.505 71.040 221.715 ;
        RECT 71.320 221.685 71.675 222.055 ;
        RECT 71.445 221.675 71.615 221.685 ;
        RECT 73.430 221.580 73.770 222.410 ;
        RECT 77.385 222.225 77.675 222.955 ;
        RECT 70.445 220.575 70.700 221.480 ;
        RECT 70.870 221.335 71.585 221.505 ;
        RECT 70.870 220.405 71.200 221.165 ;
        RECT 71.415 220.575 71.585 221.335 ;
        RECT 75.250 220.840 75.600 222.090 ;
        RECT 77.375 221.715 77.675 222.045 ;
        RECT 77.855 222.025 78.085 222.665 ;
        RECT 78.265 222.405 78.575 222.775 ;
        RECT 78.755 222.585 79.425 222.955 ;
        RECT 78.265 222.205 79.495 222.405 ;
        RECT 77.855 221.715 78.380 222.025 ;
        RECT 78.560 221.715 79.025 222.025 ;
        RECT 79.205 221.535 79.495 222.205 ;
        RECT 77.385 221.295 78.545 221.535 ;
        RECT 71.845 220.405 77.190 220.840 ;
        RECT 77.385 220.585 77.645 221.295 ;
        RECT 77.815 220.405 78.145 221.115 ;
        RECT 78.315 220.585 78.545 221.295 ;
        RECT 78.725 221.315 79.495 221.535 ;
        RECT 78.725 220.585 78.995 221.315 ;
        RECT 79.175 220.405 79.515 221.135 ;
        RECT 79.685 220.585 79.945 222.775 ;
        RECT 80.125 222.230 80.415 222.955 ;
        RECT 81.510 222.135 81.785 222.955 ;
        RECT 81.955 222.315 82.285 222.785 ;
        RECT 82.455 222.485 82.625 222.955 ;
        RECT 82.795 222.315 83.125 222.785 ;
        RECT 83.295 222.485 83.465 222.955 ;
        RECT 83.635 222.315 83.965 222.785 ;
        RECT 84.135 222.485 84.305 222.955 ;
        RECT 84.475 222.315 84.805 222.785 ;
        RECT 84.975 222.485 85.260 222.955 ;
        RECT 81.955 222.135 85.475 222.315 ;
        RECT 81.560 221.765 83.220 221.965 ;
        RECT 83.540 221.765 84.905 221.965 ;
        RECT 85.075 221.595 85.475 222.135 ;
        RECT 85.645 222.205 86.855 222.955 ;
        RECT 87.140 222.325 87.425 222.785 ;
        RECT 87.595 222.495 87.865 222.955 ;
        RECT 85.645 221.665 86.165 222.205 ;
        RECT 87.140 222.155 88.095 222.325 ;
        RECT 80.125 220.405 80.415 221.570 ;
        RECT 81.510 221.375 83.545 221.585 ;
        RECT 81.510 220.575 81.785 221.375 ;
        RECT 81.955 220.405 82.285 221.205 ;
        RECT 82.455 220.575 82.625 221.375 ;
        RECT 82.795 220.405 83.045 221.205 ;
        RECT 83.215 220.745 83.545 221.375 ;
        RECT 83.715 221.295 85.475 221.595 ;
        RECT 86.335 221.495 86.855 222.035 ;
        RECT 83.715 220.915 83.885 221.295 ;
        RECT 84.055 220.745 84.385 221.105 ;
        RECT 84.555 220.915 84.725 221.295 ;
        RECT 84.895 220.745 85.310 221.125 ;
        RECT 83.215 220.575 85.310 220.745 ;
        RECT 85.645 220.405 86.855 221.495 ;
        RECT 87.025 221.425 87.715 221.985 ;
        RECT 87.885 221.255 88.095 222.155 ;
        RECT 87.140 221.035 88.095 221.255 ;
        RECT 88.265 221.985 88.665 222.785 ;
        RECT 88.855 222.325 89.135 222.785 ;
        RECT 89.655 222.495 89.980 222.955 ;
        RECT 88.855 222.155 89.980 222.325 ;
        RECT 90.150 222.215 90.535 222.785 ;
        RECT 89.530 222.045 89.980 222.155 ;
        RECT 88.265 221.425 89.360 221.985 ;
        RECT 89.530 221.715 90.085 222.045 ;
        RECT 87.140 220.575 87.425 221.035 ;
        RECT 87.595 220.405 87.865 220.865 ;
        RECT 88.265 220.575 88.665 221.425 ;
        RECT 89.530 221.255 89.980 221.715 ;
        RECT 90.255 221.545 90.535 222.215 ;
        RECT 90.705 222.185 92.375 222.955 ;
        RECT 93.005 222.230 93.295 222.955 ;
        RECT 90.705 221.665 91.455 222.185 ;
        RECT 88.855 221.035 89.980 221.255 ;
        RECT 88.855 220.575 89.135 221.035 ;
        RECT 89.655 220.405 89.980 220.865 ;
        RECT 90.150 220.575 90.535 221.545 ;
        RECT 91.625 221.495 92.375 222.015 ;
        RECT 90.705 220.405 92.375 221.495 ;
        RECT 93.005 220.405 93.295 221.570 ;
        RECT 93.475 220.585 93.735 222.775 ;
        RECT 93.995 222.585 94.665 222.955 ;
        RECT 94.845 222.405 95.155 222.775 ;
        RECT 93.925 222.205 95.155 222.405 ;
        RECT 93.925 221.535 94.215 222.205 ;
        RECT 95.335 222.025 95.565 222.665 ;
        RECT 95.745 222.225 96.035 222.955 ;
        RECT 96.265 222.135 96.495 222.955 ;
        RECT 96.665 222.155 96.995 222.785 ;
        RECT 94.395 221.715 94.860 222.025 ;
        RECT 95.040 221.715 95.565 222.025 ;
        RECT 95.745 221.715 96.045 222.045 ;
        RECT 96.245 221.715 96.575 221.965 ;
        RECT 96.745 221.555 96.995 222.155 ;
        RECT 97.165 222.135 97.375 222.955 ;
        RECT 97.605 222.410 102.950 222.955 ;
        RECT 99.190 221.580 99.530 222.410 ;
        RECT 103.125 222.185 105.715 222.955 ;
        RECT 105.885 222.230 106.175 222.955 ;
        RECT 106.345 222.215 106.730 222.785 ;
        RECT 106.900 222.495 107.225 222.955 ;
        RECT 107.745 222.325 108.025 222.785 ;
        RECT 93.925 221.315 94.695 221.535 ;
        RECT 93.905 220.405 94.245 221.135 ;
        RECT 94.425 220.585 94.695 221.315 ;
        RECT 94.875 221.295 96.035 221.535 ;
        RECT 94.875 220.585 95.105 221.295 ;
        RECT 95.275 220.405 95.605 221.115 ;
        RECT 95.775 220.585 96.035 221.295 ;
        RECT 96.265 220.405 96.495 221.545 ;
        RECT 96.665 220.575 96.995 221.555 ;
        RECT 97.165 220.405 97.375 221.545 ;
        RECT 101.010 220.840 101.360 222.090 ;
        RECT 103.125 221.665 104.335 222.185 ;
        RECT 104.505 221.495 105.715 222.015 ;
        RECT 97.605 220.405 102.950 220.840 ;
        RECT 103.125 220.405 105.715 221.495 ;
        RECT 105.885 220.405 106.175 221.570 ;
        RECT 106.345 221.545 106.625 222.215 ;
        RECT 106.900 222.155 108.025 222.325 ;
        RECT 106.900 222.045 107.350 222.155 ;
        RECT 106.795 221.715 107.350 222.045 ;
        RECT 108.215 221.985 108.615 222.785 ;
        RECT 109.015 222.495 109.285 222.955 ;
        RECT 109.455 222.325 109.740 222.785 ;
        RECT 106.345 220.575 106.730 221.545 ;
        RECT 106.900 221.255 107.350 221.715 ;
        RECT 107.520 221.425 108.615 221.985 ;
        RECT 106.900 221.035 108.025 221.255 ;
        RECT 106.900 220.405 107.225 220.865 ;
        RECT 107.745 220.575 108.025 221.035 ;
        RECT 108.215 220.575 108.615 221.425 ;
        RECT 108.785 222.155 109.740 222.325 ;
        RECT 108.785 221.255 108.995 222.155 ;
        RECT 110.065 222.135 110.295 222.955 ;
        RECT 110.465 222.155 110.795 222.785 ;
        RECT 109.165 221.425 109.855 221.985 ;
        RECT 110.045 221.715 110.375 221.965 ;
        RECT 110.545 221.555 110.795 222.155 ;
        RECT 110.965 222.135 111.175 222.955 ;
        RECT 111.405 222.185 113.075 222.955 ;
        RECT 111.405 221.665 112.155 222.185 ;
        RECT 108.785 221.035 109.740 221.255 ;
        RECT 109.015 220.405 109.285 220.865 ;
        RECT 109.455 220.575 109.740 221.035 ;
        RECT 110.065 220.405 110.295 221.545 ;
        RECT 110.465 220.575 110.795 221.555 ;
        RECT 110.965 220.405 111.175 221.545 ;
        RECT 112.325 221.495 113.075 222.015 ;
        RECT 111.405 220.405 113.075 221.495 ;
        RECT 113.725 221.375 113.955 222.715 ;
        RECT 114.135 221.875 114.365 222.775 ;
        RECT 114.565 222.175 114.810 222.955 ;
        RECT 114.980 222.415 115.410 222.775 ;
        RECT 115.990 222.585 116.720 222.955 ;
        RECT 114.980 222.225 116.720 222.415 ;
        RECT 114.980 221.995 115.200 222.225 ;
        RECT 114.135 221.195 114.475 221.875 ;
        RECT 113.725 220.995 114.475 221.195 ;
        RECT 114.655 221.695 115.200 221.995 ;
        RECT 113.725 220.605 113.965 220.995 ;
        RECT 114.135 220.405 114.485 220.815 ;
        RECT 114.655 220.585 114.985 221.695 ;
        RECT 115.370 221.425 115.795 222.045 ;
        RECT 115.990 221.425 116.250 222.045 ;
        RECT 116.460 221.715 116.720 222.225 ;
        RECT 115.155 221.055 116.180 221.255 ;
        RECT 115.155 220.585 115.335 221.055 ;
        RECT 115.505 220.405 115.835 220.885 ;
        RECT 116.010 220.585 116.180 221.055 ;
        RECT 116.445 220.405 116.730 221.545 ;
        RECT 116.920 220.585 117.200 222.775 ;
        RECT 117.385 222.205 118.595 222.955 ;
        RECT 118.765 222.230 119.055 222.955 ;
        RECT 117.385 221.665 117.905 222.205 ;
        RECT 119.225 222.185 122.735 222.955 ;
        RECT 123.105 222.325 123.435 222.685 ;
        RECT 124.055 222.495 124.305 222.955 ;
        RECT 124.475 222.495 125.035 222.785 ;
        RECT 118.075 221.495 118.595 222.035 ;
        RECT 119.225 221.665 120.875 222.185 ;
        RECT 123.105 222.135 124.495 222.325 ;
        RECT 124.325 222.045 124.495 222.135 ;
        RECT 117.385 220.405 118.595 221.495 ;
        RECT 118.765 220.405 119.055 221.570 ;
        RECT 121.045 221.495 122.735 222.015 ;
        RECT 119.225 220.405 122.735 221.495 ;
        RECT 122.920 221.715 123.595 221.965 ;
        RECT 123.815 221.715 124.155 221.965 ;
        RECT 124.325 221.715 124.615 222.045 ;
        RECT 122.920 221.355 123.185 221.715 ;
        RECT 123.885 221.675 124.055 221.715 ;
        RECT 124.325 221.465 124.495 221.715 ;
        RECT 122.965 221.335 123.135 221.355 ;
        RECT 123.555 221.295 124.495 221.465 ;
        RECT 123.105 220.405 123.385 221.075 ;
        RECT 123.555 220.745 123.855 221.295 ;
        RECT 124.785 221.125 125.035 222.495 ;
        RECT 124.055 220.405 124.385 221.125 ;
        RECT 124.575 220.575 125.035 221.125 ;
        RECT 125.205 222.280 125.465 222.785 ;
        RECT 125.645 222.575 125.975 222.955 ;
        RECT 126.155 222.405 126.325 222.785 ;
        RECT 125.205 221.480 125.375 222.280 ;
        RECT 125.660 222.235 126.325 222.405 ;
        RECT 126.585 222.280 126.845 222.785 ;
        RECT 127.025 222.575 127.355 222.955 ;
        RECT 127.535 222.405 127.705 222.785 ;
        RECT 125.660 221.980 125.830 222.235 ;
        RECT 125.545 221.650 125.830 221.980 ;
        RECT 126.065 221.685 126.395 222.055 ;
        RECT 126.185 221.675 126.355 221.685 ;
        RECT 125.660 221.505 125.830 221.650 ;
        RECT 126.585 221.505 126.755 222.280 ;
        RECT 127.040 222.235 127.705 222.405 ;
        RECT 127.040 221.980 127.210 222.235 ;
        RECT 127.965 222.185 131.475 222.955 ;
        RECT 131.645 222.230 131.935 222.955 ;
        RECT 133.025 222.280 133.285 222.785 ;
        RECT 133.465 222.575 133.795 222.955 ;
        RECT 133.975 222.405 134.145 222.785 ;
        RECT 126.925 221.650 127.210 221.980 ;
        RECT 127.445 221.685 127.775 222.055 ;
        RECT 127.565 221.675 127.735 221.685 ;
        RECT 127.965 221.665 129.615 222.185 ;
        RECT 127.040 221.505 127.210 221.650 ;
        RECT 125.205 220.575 125.475 221.480 ;
        RECT 125.660 221.335 126.325 221.505 ;
        RECT 125.645 220.405 125.975 221.165 ;
        RECT 126.155 220.575 126.325 221.335 ;
        RECT 126.585 221.480 126.815 221.505 ;
        RECT 126.585 220.575 126.855 221.480 ;
        RECT 127.040 221.335 127.705 221.505 ;
        RECT 129.785 221.495 131.475 222.015 ;
        RECT 127.025 220.405 127.355 221.165 ;
        RECT 127.535 220.575 127.705 221.335 ;
        RECT 127.965 220.405 131.475 221.495 ;
        RECT 131.645 220.405 131.935 221.570 ;
        RECT 133.025 221.480 133.195 222.280 ;
        RECT 133.480 222.235 134.145 222.405 ;
        RECT 133.480 221.980 133.650 222.235 ;
        RECT 134.410 222.215 134.665 222.785 ;
        RECT 134.835 222.555 135.165 222.955 ;
        RECT 135.590 222.420 136.120 222.785 ;
        RECT 135.590 222.385 135.765 222.420 ;
        RECT 134.835 222.215 135.765 222.385 ;
        RECT 133.365 221.650 133.650 221.980 ;
        RECT 133.885 221.685 134.215 222.055 ;
        RECT 134.005 221.675 134.175 221.685 ;
        RECT 133.480 221.505 133.650 221.650 ;
        RECT 134.410 221.545 134.580 222.215 ;
        RECT 134.835 222.045 135.005 222.215 ;
        RECT 134.750 221.715 135.005 222.045 ;
        RECT 135.230 221.715 135.425 222.045 ;
        RECT 133.025 220.575 133.295 221.480 ;
        RECT 133.480 221.335 134.145 221.505 ;
        RECT 133.465 220.405 133.795 221.165 ;
        RECT 133.975 220.575 134.145 221.335 ;
        RECT 134.410 220.575 134.745 221.545 ;
        RECT 134.915 220.405 135.085 221.545 ;
        RECT 135.255 220.745 135.425 221.715 ;
        RECT 135.595 221.085 135.765 222.215 ;
        RECT 135.935 221.425 136.105 222.225 ;
        RECT 136.310 221.845 136.585 222.785 ;
        RECT 136.305 221.675 136.585 221.845 ;
        RECT 136.310 221.625 136.585 221.675 ;
        RECT 136.755 221.425 136.945 222.785 ;
        RECT 137.125 222.420 137.635 222.955 ;
        RECT 137.855 222.145 138.100 222.750 ;
        RECT 138.545 222.215 138.930 222.785 ;
        RECT 139.100 222.495 139.425 222.955 ;
        RECT 139.945 222.325 140.225 222.785 ;
        RECT 137.145 221.975 138.375 222.145 ;
        RECT 135.935 221.255 136.945 221.425 ;
        RECT 137.115 221.410 137.865 221.600 ;
        RECT 137.115 221.335 137.395 221.410 ;
        RECT 135.595 220.915 136.720 221.085 ;
        RECT 137.115 220.745 137.285 221.335 ;
        RECT 138.035 221.165 138.375 221.975 ;
        RECT 135.255 220.575 137.285 220.745 ;
        RECT 137.455 220.405 137.625 221.165 ;
        RECT 137.860 220.755 138.375 221.165 ;
        RECT 138.545 221.545 138.825 222.215 ;
        RECT 139.100 222.155 140.225 222.325 ;
        RECT 139.100 222.045 139.550 222.155 ;
        RECT 138.995 221.715 139.550 222.045 ;
        RECT 140.415 221.985 140.815 222.785 ;
        RECT 141.215 222.495 141.485 222.955 ;
        RECT 141.655 222.325 141.940 222.785 ;
        RECT 138.545 220.575 138.930 221.545 ;
        RECT 139.100 221.255 139.550 221.715 ;
        RECT 139.720 221.425 140.815 221.985 ;
        RECT 139.100 221.035 140.225 221.255 ;
        RECT 139.100 220.405 139.425 220.865 ;
        RECT 139.945 220.575 140.225 221.035 ;
        RECT 140.415 220.575 140.815 221.425 ;
        RECT 140.985 222.155 141.940 222.325 ;
        RECT 142.225 222.280 142.485 222.785 ;
        RECT 142.665 222.575 142.995 222.955 ;
        RECT 143.175 222.405 143.345 222.785 ;
        RECT 140.985 221.255 141.195 222.155 ;
        RECT 141.365 221.425 142.055 221.985 ;
        RECT 142.225 221.480 142.395 222.280 ;
        RECT 142.680 222.235 143.345 222.405 ;
        RECT 142.680 221.980 142.850 222.235 ;
        RECT 144.525 222.230 144.815 222.955 ;
        RECT 145.260 222.145 145.505 222.750 ;
        RECT 145.725 222.420 146.235 222.955 ;
        RECT 142.565 221.650 142.850 221.980 ;
        RECT 143.085 221.685 143.415 222.055 ;
        RECT 144.985 221.975 146.215 222.145 ;
        RECT 143.205 221.675 143.375 221.685 ;
        RECT 142.680 221.505 142.850 221.650 ;
        RECT 140.985 221.035 141.940 221.255 ;
        RECT 141.215 220.405 141.485 220.865 ;
        RECT 141.655 220.575 141.940 221.035 ;
        RECT 142.225 220.575 142.495 221.480 ;
        RECT 142.680 221.335 143.345 221.505 ;
        RECT 142.665 220.405 142.995 221.165 ;
        RECT 143.175 220.575 143.345 221.335 ;
        RECT 144.525 220.405 144.815 221.570 ;
        RECT 144.985 221.165 145.325 221.975 ;
        RECT 145.495 221.410 146.245 221.600 ;
        RECT 145.505 221.335 145.675 221.410 ;
        RECT 144.985 220.755 145.500 221.165 ;
        RECT 145.735 220.405 145.905 221.165 ;
        RECT 146.075 220.745 146.245 221.410 ;
        RECT 146.415 221.425 146.605 222.785 ;
        RECT 146.775 222.185 147.050 222.785 ;
        RECT 147.240 222.420 147.770 222.785 ;
        RECT 148.195 222.555 148.525 222.955 ;
        RECT 147.595 222.385 147.770 222.420 ;
        RECT 146.775 222.015 147.055 222.185 ;
        RECT 146.775 221.625 147.050 222.015 ;
        RECT 147.255 221.425 147.425 222.225 ;
        RECT 146.415 221.255 147.425 221.425 ;
        RECT 147.595 222.215 148.525 222.385 ;
        RECT 148.695 222.215 148.950 222.785 ;
        RECT 147.595 221.085 147.765 222.215 ;
        RECT 148.355 222.045 148.525 222.215 ;
        RECT 146.640 220.915 147.765 221.085 ;
        RECT 147.935 221.715 148.130 222.045 ;
        RECT 148.355 221.715 148.610 222.045 ;
        RECT 147.935 220.745 148.105 221.715 ;
        RECT 148.780 221.545 148.950 222.215 ;
        RECT 149.400 222.145 149.645 222.750 ;
        RECT 149.865 222.420 150.375 222.955 ;
        RECT 146.075 220.575 148.105 220.745 ;
        RECT 148.275 220.405 148.445 221.545 ;
        RECT 148.615 220.575 148.950 221.545 ;
        RECT 149.125 221.975 150.355 222.145 ;
        RECT 149.125 221.165 149.465 221.975 ;
        RECT 149.635 221.410 150.385 221.600 ;
        RECT 149.645 221.335 149.815 221.410 ;
        RECT 149.125 220.755 149.640 221.165 ;
        RECT 149.875 220.405 150.045 221.165 ;
        RECT 150.215 220.745 150.385 221.410 ;
        RECT 150.555 221.425 150.745 222.785 ;
        RECT 150.915 221.845 151.190 222.785 ;
        RECT 151.380 222.420 151.910 222.785 ;
        RECT 152.335 222.555 152.665 222.955 ;
        RECT 151.735 222.385 151.910 222.420 ;
        RECT 150.915 221.675 151.195 221.845 ;
        RECT 150.915 221.625 151.190 221.675 ;
        RECT 151.395 221.425 151.565 222.225 ;
        RECT 150.555 221.255 151.565 221.425 ;
        RECT 151.735 222.215 152.665 222.385 ;
        RECT 152.835 222.215 153.090 222.785 ;
        RECT 151.735 221.085 151.905 222.215 ;
        RECT 152.495 222.045 152.665 222.215 ;
        RECT 150.780 220.915 151.905 221.085 ;
        RECT 152.075 221.715 152.270 222.045 ;
        RECT 152.495 221.715 152.750 222.045 ;
        RECT 152.075 220.745 152.245 221.715 ;
        RECT 152.920 221.545 153.090 222.215 ;
        RECT 150.215 220.575 152.245 220.745 ;
        RECT 152.415 220.405 152.585 221.545 ;
        RECT 152.755 220.575 153.090 221.545 ;
        RECT 153.265 222.215 153.650 222.785 ;
        RECT 153.820 222.495 154.145 222.955 ;
        RECT 154.665 222.325 154.945 222.785 ;
        RECT 153.265 221.545 153.545 222.215 ;
        RECT 153.820 222.155 154.945 222.325 ;
        RECT 153.820 222.045 154.270 222.155 ;
        RECT 153.715 221.715 154.270 222.045 ;
        RECT 155.135 221.985 155.535 222.785 ;
        RECT 155.935 222.495 156.205 222.955 ;
        RECT 156.375 222.325 156.660 222.785 ;
        RECT 153.265 220.575 153.650 221.545 ;
        RECT 153.820 221.255 154.270 221.715 ;
        RECT 154.440 221.425 155.535 221.985 ;
        RECT 153.820 221.035 154.945 221.255 ;
        RECT 153.820 220.405 154.145 220.865 ;
        RECT 154.665 220.575 154.945 221.035 ;
        RECT 155.135 220.575 155.535 221.425 ;
        RECT 155.705 222.155 156.660 222.325 ;
        RECT 156.945 222.205 158.155 222.955 ;
        RECT 155.705 221.255 155.915 222.155 ;
        RECT 156.085 221.425 156.775 221.985 ;
        RECT 156.945 221.495 157.465 222.035 ;
        RECT 157.635 221.665 158.155 222.205 ;
        RECT 155.705 221.035 156.660 221.255 ;
        RECT 155.935 220.405 156.205 220.865 ;
        RECT 156.375 220.575 156.660 221.035 ;
        RECT 156.945 220.405 158.155 221.495 ;
        RECT 2.760 220.235 158.240 220.405 ;
        RECT 2.845 219.145 4.055 220.235 ;
        RECT 4.225 219.800 9.570 220.235 ;
        RECT 9.745 219.800 15.090 220.235 ;
        RECT 2.845 218.435 3.365 218.975 ;
        RECT 3.535 218.605 4.055 219.145 ;
        RECT 2.845 217.685 4.055 218.435 ;
        RECT 5.810 218.230 6.150 219.060 ;
        RECT 7.630 218.550 7.980 219.800 ;
        RECT 11.330 218.230 11.670 219.060 ;
        RECT 13.150 218.550 13.500 219.800 ;
        RECT 15.725 219.070 16.015 220.235 ;
        RECT 16.185 219.800 21.530 220.235 ;
        RECT 21.705 219.800 27.050 220.235 ;
        RECT 27.225 219.800 32.570 220.235 ;
        RECT 32.745 219.800 38.090 220.235 ;
        RECT 4.225 217.685 9.570 218.230 ;
        RECT 9.745 217.685 15.090 218.230 ;
        RECT 15.725 217.685 16.015 218.410 ;
        RECT 17.770 218.230 18.110 219.060 ;
        RECT 19.590 218.550 19.940 219.800 ;
        RECT 23.290 218.230 23.630 219.060 ;
        RECT 25.110 218.550 25.460 219.800 ;
        RECT 28.810 218.230 29.150 219.060 ;
        RECT 30.630 218.550 30.980 219.800 ;
        RECT 34.330 218.230 34.670 219.060 ;
        RECT 36.150 218.550 36.500 219.800 ;
        RECT 38.265 219.145 40.855 220.235 ;
        RECT 38.265 218.455 39.475 218.975 ;
        RECT 39.645 218.625 40.855 219.145 ;
        RECT 41.485 219.070 41.775 220.235 ;
        RECT 41.945 219.800 47.290 220.235 ;
        RECT 47.465 219.800 52.810 220.235 ;
        RECT 16.185 217.685 21.530 218.230 ;
        RECT 21.705 217.685 27.050 218.230 ;
        RECT 27.225 217.685 32.570 218.230 ;
        RECT 32.745 217.685 38.090 218.230 ;
        RECT 38.265 217.685 40.855 218.455 ;
        RECT 41.485 217.685 41.775 218.410 ;
        RECT 43.530 218.230 43.870 219.060 ;
        RECT 45.350 218.550 45.700 219.800 ;
        RECT 49.050 218.230 49.390 219.060 ;
        RECT 50.870 218.550 51.220 219.800 ;
        RECT 52.985 219.145 54.195 220.235 ;
        RECT 52.985 218.435 53.505 218.975 ;
        RECT 53.675 218.605 54.195 219.145 ;
        RECT 54.405 219.095 54.635 220.235 ;
        RECT 54.805 219.085 55.135 220.065 ;
        RECT 55.305 219.095 55.515 220.235 ;
        RECT 55.800 219.365 56.085 220.235 ;
        RECT 56.255 219.605 56.515 220.065 ;
        RECT 56.690 219.775 56.945 220.235 ;
        RECT 57.115 219.605 57.375 220.065 ;
        RECT 56.255 219.435 57.375 219.605 ;
        RECT 57.545 219.435 57.855 220.235 ;
        RECT 56.255 219.185 56.515 219.435 ;
        RECT 58.025 219.265 58.335 220.065 ;
        RECT 58.595 219.565 58.765 220.065 ;
        RECT 58.935 219.735 59.265 220.235 ;
        RECT 58.595 219.395 59.260 219.565 ;
        RECT 54.385 218.675 54.715 218.925 ;
        RECT 41.945 217.685 47.290 218.230 ;
        RECT 47.465 217.685 52.810 218.230 ;
        RECT 52.985 217.685 54.195 218.435 ;
        RECT 54.405 217.685 54.635 218.505 ;
        RECT 54.885 218.485 55.135 219.085 ;
        RECT 55.760 219.015 56.515 219.185 ;
        RECT 57.305 219.095 58.335 219.265 ;
        RECT 55.760 218.505 56.165 219.015 ;
        RECT 57.305 218.845 57.475 219.095 ;
        RECT 56.335 218.675 57.475 218.845 ;
        RECT 54.805 217.855 55.135 218.485 ;
        RECT 55.305 217.685 55.515 218.505 ;
        RECT 55.760 218.335 57.410 218.505 ;
        RECT 57.645 218.355 57.995 218.925 ;
        RECT 55.805 217.685 56.085 218.165 ;
        RECT 56.255 217.945 56.515 218.335 ;
        RECT 56.690 217.685 56.945 218.165 ;
        RECT 57.115 217.945 57.410 218.335 ;
        RECT 58.165 218.185 58.335 219.095 ;
        RECT 58.510 218.575 58.860 219.225 ;
        RECT 59.030 218.405 59.260 219.395 ;
        RECT 57.590 217.685 57.865 218.165 ;
        RECT 58.035 217.855 58.335 218.185 ;
        RECT 58.595 218.235 59.260 218.405 ;
        RECT 58.595 217.945 58.765 218.235 ;
        RECT 58.935 217.685 59.265 218.065 ;
        RECT 59.435 217.945 59.620 220.065 ;
        RECT 59.860 219.775 60.125 220.235 ;
        RECT 60.295 219.640 60.545 220.065 ;
        RECT 60.755 219.790 61.860 219.960 ;
        RECT 60.240 219.510 60.545 219.640 ;
        RECT 59.790 218.315 60.070 219.265 ;
        RECT 60.240 218.405 60.410 219.510 ;
        RECT 60.580 218.725 60.820 219.320 ;
        RECT 60.990 219.255 61.520 219.620 ;
        RECT 60.990 218.555 61.160 219.255 ;
        RECT 61.690 219.175 61.860 219.790 ;
        RECT 62.030 219.435 62.200 220.235 ;
        RECT 62.370 219.735 62.620 220.065 ;
        RECT 62.845 219.765 63.730 219.935 ;
        RECT 61.690 219.085 62.200 219.175 ;
        RECT 60.240 218.275 60.465 218.405 ;
        RECT 60.635 218.335 61.160 218.555 ;
        RECT 61.330 218.915 62.200 219.085 ;
        RECT 59.875 217.685 60.125 218.145 ;
        RECT 60.295 218.135 60.465 218.275 ;
        RECT 61.330 218.135 61.500 218.915 ;
        RECT 62.030 218.845 62.200 218.915 ;
        RECT 61.710 218.665 61.910 218.695 ;
        RECT 62.370 218.665 62.540 219.735 ;
        RECT 62.710 218.845 62.900 219.565 ;
        RECT 61.710 218.365 62.540 218.665 ;
        RECT 63.070 218.635 63.390 219.595 ;
        RECT 60.295 217.965 60.630 218.135 ;
        RECT 60.825 217.965 61.500 218.135 ;
        RECT 61.820 217.685 62.190 218.185 ;
        RECT 62.370 218.135 62.540 218.365 ;
        RECT 62.925 218.305 63.390 218.635 ;
        RECT 63.560 218.925 63.730 219.765 ;
        RECT 63.910 219.735 64.225 220.235 ;
        RECT 64.455 219.505 64.795 220.065 ;
        RECT 63.900 219.130 64.795 219.505 ;
        RECT 64.965 219.225 65.135 220.235 ;
        RECT 64.605 218.925 64.795 219.130 ;
        RECT 65.305 219.175 65.635 220.020 ;
        RECT 65.305 219.095 65.695 219.175 ;
        RECT 65.865 219.145 67.075 220.235 ;
        RECT 65.480 219.045 65.695 219.095 ;
        RECT 63.560 218.595 64.435 218.925 ;
        RECT 64.605 218.595 65.355 218.925 ;
        RECT 63.560 218.135 63.730 218.595 ;
        RECT 64.605 218.425 64.805 218.595 ;
        RECT 65.525 218.465 65.695 219.045 ;
        RECT 65.470 218.445 65.695 218.465 ;
        RECT 65.465 218.425 65.695 218.445 ;
        RECT 62.370 217.965 62.775 218.135 ;
        RECT 62.945 217.965 63.730 218.135 ;
        RECT 64.005 217.685 64.215 218.215 ;
        RECT 64.475 217.900 64.805 218.425 ;
        RECT 65.315 218.340 65.695 218.425 ;
        RECT 65.865 218.435 66.385 218.975 ;
        RECT 66.555 218.605 67.075 219.145 ;
        RECT 67.245 219.070 67.535 220.235 ;
        RECT 67.760 219.365 68.045 220.235 ;
        RECT 68.215 219.605 68.475 220.065 ;
        RECT 68.650 219.775 68.905 220.235 ;
        RECT 69.075 219.605 69.335 220.065 ;
        RECT 68.215 219.435 69.335 219.605 ;
        RECT 69.505 219.435 69.815 220.235 ;
        RECT 68.215 219.185 68.475 219.435 ;
        RECT 69.985 219.265 70.295 220.065 ;
        RECT 70.630 219.895 72.725 220.065 ;
        RECT 70.630 219.515 71.045 219.895 ;
        RECT 71.215 219.345 71.385 219.725 ;
        RECT 71.555 219.535 71.885 219.895 ;
        RECT 72.055 219.345 72.225 219.725 ;
        RECT 67.720 219.015 68.475 219.185 ;
        RECT 69.265 219.095 70.295 219.265 ;
        RECT 67.720 218.505 68.125 219.015 ;
        RECT 69.265 218.845 69.435 219.095 ;
        RECT 68.295 218.675 69.435 218.845 ;
        RECT 64.975 217.685 65.145 218.295 ;
        RECT 65.315 217.905 65.645 218.340 ;
        RECT 65.865 217.685 67.075 218.435 ;
        RECT 67.245 217.685 67.535 218.410 ;
        RECT 67.720 218.335 69.370 218.505 ;
        RECT 69.605 218.355 69.955 218.925 ;
        RECT 67.765 217.685 68.045 218.165 ;
        RECT 68.215 217.945 68.475 218.335 ;
        RECT 68.650 217.685 68.905 218.165 ;
        RECT 69.075 217.945 69.370 218.335 ;
        RECT 70.125 218.185 70.295 219.095 ;
        RECT 70.465 219.045 72.225 219.345 ;
        RECT 72.395 219.265 72.725 219.895 ;
        RECT 72.895 219.435 73.145 220.235 ;
        RECT 73.315 219.265 73.485 220.065 ;
        RECT 73.655 219.435 73.985 220.235 ;
        RECT 74.155 219.265 74.430 220.065 ;
        RECT 72.395 219.055 74.430 219.265 ;
        RECT 75.105 219.095 75.335 220.235 ;
        RECT 75.505 219.085 75.835 220.065 ;
        RECT 76.005 219.095 76.215 220.235 ;
        RECT 70.465 218.505 70.865 219.045 ;
        RECT 71.035 218.675 72.400 218.875 ;
        RECT 72.720 218.675 74.380 218.875 ;
        RECT 75.085 218.675 75.415 218.925 ;
        RECT 70.465 218.325 73.985 218.505 ;
        RECT 69.550 217.685 69.825 218.165 ;
        RECT 69.995 217.855 70.295 218.185 ;
        RECT 70.680 217.685 70.965 218.155 ;
        RECT 71.135 217.855 71.465 218.325 ;
        RECT 71.635 217.685 71.805 218.155 ;
        RECT 71.975 217.855 72.305 218.325 ;
        RECT 72.475 217.685 72.645 218.155 ;
        RECT 72.815 217.855 73.145 218.325 ;
        RECT 73.315 217.685 73.485 218.155 ;
        RECT 73.655 217.855 73.985 218.325 ;
        RECT 74.155 217.685 74.430 218.505 ;
        RECT 75.105 217.685 75.335 218.505 ;
        RECT 75.585 218.485 75.835 219.085 ;
        RECT 75.505 217.855 75.835 218.485 ;
        RECT 76.005 217.685 76.215 218.505 ;
        RECT 76.455 217.865 76.715 220.055 ;
        RECT 76.885 219.505 77.225 220.235 ;
        RECT 77.405 219.325 77.675 220.055 ;
        RECT 76.905 219.105 77.675 219.325 ;
        RECT 77.855 219.345 78.085 220.055 ;
        RECT 78.255 219.525 78.585 220.235 ;
        RECT 78.755 219.345 79.015 220.055 ;
        RECT 79.295 219.565 79.465 220.065 ;
        RECT 79.635 219.735 79.965 220.235 ;
        RECT 79.295 219.395 79.960 219.565 ;
        RECT 77.855 219.105 79.015 219.345 ;
        RECT 76.905 218.435 77.195 219.105 ;
        RECT 77.375 218.615 77.840 218.925 ;
        RECT 78.020 218.615 78.545 218.925 ;
        RECT 76.905 218.235 78.135 218.435 ;
        RECT 76.975 217.685 77.645 218.055 ;
        RECT 77.825 217.865 78.135 218.235 ;
        RECT 78.315 217.975 78.545 218.615 ;
        RECT 78.725 218.595 79.025 218.925 ;
        RECT 79.210 218.575 79.560 219.225 ;
        RECT 78.725 217.685 79.015 218.415 ;
        RECT 79.730 218.405 79.960 219.395 ;
        RECT 79.295 218.235 79.960 218.405 ;
        RECT 79.295 217.945 79.465 218.235 ;
        RECT 79.635 217.685 79.965 218.065 ;
        RECT 80.135 217.945 80.320 220.065 ;
        RECT 80.560 219.775 80.825 220.235 ;
        RECT 80.995 219.640 81.245 220.065 ;
        RECT 81.455 219.790 82.560 219.960 ;
        RECT 80.940 219.510 81.245 219.640 ;
        RECT 80.490 218.315 80.770 219.265 ;
        RECT 80.940 218.405 81.110 219.510 ;
        RECT 81.280 218.725 81.520 219.320 ;
        RECT 81.690 219.255 82.220 219.620 ;
        RECT 81.690 218.555 81.860 219.255 ;
        RECT 82.390 219.175 82.560 219.790 ;
        RECT 82.730 219.435 82.900 220.235 ;
        RECT 83.070 219.735 83.320 220.065 ;
        RECT 83.545 219.765 84.430 219.935 ;
        RECT 82.390 219.085 82.900 219.175 ;
        RECT 80.940 218.275 81.165 218.405 ;
        RECT 81.335 218.335 81.860 218.555 ;
        RECT 82.030 218.915 82.900 219.085 ;
        RECT 80.575 217.685 80.825 218.145 ;
        RECT 80.995 218.135 81.165 218.275 ;
        RECT 82.030 218.135 82.200 218.915 ;
        RECT 82.730 218.845 82.900 218.915 ;
        RECT 82.410 218.665 82.610 218.695 ;
        RECT 83.070 218.665 83.240 219.735 ;
        RECT 83.410 218.845 83.600 219.565 ;
        RECT 82.410 218.365 83.240 218.665 ;
        RECT 83.770 218.635 84.090 219.595 ;
        RECT 80.995 217.965 81.330 218.135 ;
        RECT 81.525 217.965 82.200 218.135 ;
        RECT 82.520 217.685 82.890 218.185 ;
        RECT 83.070 218.135 83.240 218.365 ;
        RECT 83.625 218.305 84.090 218.635 ;
        RECT 84.260 218.925 84.430 219.765 ;
        RECT 84.610 219.735 84.925 220.235 ;
        RECT 85.155 219.505 85.495 220.065 ;
        RECT 84.600 219.130 85.495 219.505 ;
        RECT 85.665 219.225 85.835 220.235 ;
        RECT 85.305 218.925 85.495 219.130 ;
        RECT 86.005 219.175 86.335 220.020 ;
        RECT 86.505 219.320 86.675 220.235 ;
        RECT 87.190 219.895 89.285 220.065 ;
        RECT 87.190 219.515 87.605 219.895 ;
        RECT 87.775 219.345 87.945 219.725 ;
        RECT 88.115 219.535 88.445 219.895 ;
        RECT 88.615 219.345 88.785 219.725 ;
        RECT 86.005 219.095 86.395 219.175 ;
        RECT 86.180 219.045 86.395 219.095 ;
        RECT 84.260 218.595 85.135 218.925 ;
        RECT 85.305 218.595 86.055 218.925 ;
        RECT 84.260 218.135 84.430 218.595 ;
        RECT 85.305 218.425 85.505 218.595 ;
        RECT 86.225 218.465 86.395 219.045 ;
        RECT 86.170 218.425 86.395 218.465 ;
        RECT 83.070 217.965 83.475 218.135 ;
        RECT 83.645 217.965 84.430 218.135 ;
        RECT 84.705 217.685 84.915 218.215 ;
        RECT 85.175 217.900 85.505 218.425 ;
        RECT 86.015 218.340 86.395 218.425 ;
        RECT 87.025 219.045 88.785 219.345 ;
        RECT 88.955 219.265 89.285 219.895 ;
        RECT 89.455 219.435 89.705 220.235 ;
        RECT 89.875 219.265 90.045 220.065 ;
        RECT 90.215 219.435 90.545 220.235 ;
        RECT 90.715 219.265 90.990 220.065 ;
        RECT 88.955 219.055 90.990 219.265 ;
        RECT 91.165 219.145 92.835 220.235 ;
        RECT 87.025 218.505 87.425 219.045 ;
        RECT 87.595 218.675 88.960 218.875 ;
        RECT 89.280 218.675 90.940 218.875 ;
        RECT 85.675 217.685 85.845 218.295 ;
        RECT 86.015 217.905 86.345 218.340 ;
        RECT 87.025 218.325 90.545 218.505 ;
        RECT 86.515 217.685 86.685 218.200 ;
        RECT 87.240 217.685 87.525 218.155 ;
        RECT 87.695 217.855 88.025 218.325 ;
        RECT 88.195 217.685 88.365 218.155 ;
        RECT 88.535 217.855 88.865 218.325 ;
        RECT 89.035 217.685 89.205 218.155 ;
        RECT 89.375 217.855 89.705 218.325 ;
        RECT 89.875 217.685 90.045 218.155 ;
        RECT 90.215 217.855 90.545 218.325 ;
        RECT 90.715 217.685 90.990 218.505 ;
        RECT 91.165 218.455 91.915 218.975 ;
        RECT 92.085 218.625 92.835 219.145 ;
        RECT 93.005 219.070 93.295 220.235 ;
        RECT 93.580 219.605 93.865 220.065 ;
        RECT 94.035 219.775 94.305 220.235 ;
        RECT 93.580 219.385 94.535 219.605 ;
        RECT 93.465 218.655 94.155 219.215 ;
        RECT 94.325 218.485 94.535 219.385 ;
        RECT 91.165 217.685 92.835 218.455 ;
        RECT 93.005 217.685 93.295 218.410 ;
        RECT 93.580 218.315 94.535 218.485 ;
        RECT 94.705 219.215 95.105 220.065 ;
        RECT 95.295 219.605 95.575 220.065 ;
        RECT 96.095 219.775 96.420 220.235 ;
        RECT 95.295 219.385 96.420 219.605 ;
        RECT 94.705 218.655 95.800 219.215 ;
        RECT 95.970 218.925 96.420 219.385 ;
        RECT 96.590 219.095 96.975 220.065 ;
        RECT 93.580 217.855 93.865 218.315 ;
        RECT 94.035 217.685 94.305 218.145 ;
        RECT 94.705 217.855 95.105 218.655 ;
        RECT 95.970 218.595 96.525 218.925 ;
        RECT 95.970 218.485 96.420 218.595 ;
        RECT 95.295 218.315 96.420 218.485 ;
        RECT 96.695 218.425 96.975 219.095 ;
        RECT 95.295 217.855 95.575 218.315 ;
        RECT 96.095 217.685 96.420 218.145 ;
        RECT 96.590 217.855 96.975 218.425 ;
        RECT 97.155 217.865 97.415 220.055 ;
        RECT 97.585 219.505 97.925 220.235 ;
        RECT 98.105 219.325 98.375 220.055 ;
        RECT 97.605 219.105 98.375 219.325 ;
        RECT 98.555 219.345 98.785 220.055 ;
        RECT 98.955 219.525 99.285 220.235 ;
        RECT 99.455 219.345 99.715 220.055 ;
        RECT 100.455 219.565 100.625 220.065 ;
        RECT 100.795 219.735 101.125 220.235 ;
        RECT 100.455 219.395 101.120 219.565 ;
        RECT 98.555 219.105 99.715 219.345 ;
        RECT 97.605 218.435 97.895 219.105 ;
        RECT 98.075 218.615 98.540 218.925 ;
        RECT 98.720 218.615 99.245 218.925 ;
        RECT 97.605 218.235 98.835 218.435 ;
        RECT 97.675 217.685 98.345 218.055 ;
        RECT 98.525 217.865 98.835 218.235 ;
        RECT 99.015 217.975 99.245 218.615 ;
        RECT 99.425 218.595 99.725 218.925 ;
        RECT 100.370 218.575 100.720 219.225 ;
        RECT 99.425 217.685 99.715 218.415 ;
        RECT 100.890 218.405 101.120 219.395 ;
        RECT 100.455 218.235 101.120 218.405 ;
        RECT 100.455 217.945 100.625 218.235 ;
        RECT 100.795 217.685 101.125 218.065 ;
        RECT 101.295 217.945 101.480 220.065 ;
        RECT 101.720 219.775 101.985 220.235 ;
        RECT 102.155 219.640 102.405 220.065 ;
        RECT 102.615 219.790 103.720 219.960 ;
        RECT 102.100 219.510 102.405 219.640 ;
        RECT 101.650 218.315 101.930 219.265 ;
        RECT 102.100 218.405 102.270 219.510 ;
        RECT 102.440 218.725 102.680 219.320 ;
        RECT 102.850 219.255 103.380 219.620 ;
        RECT 102.850 218.555 103.020 219.255 ;
        RECT 103.550 219.175 103.720 219.790 ;
        RECT 103.890 219.435 104.060 220.235 ;
        RECT 104.230 219.735 104.480 220.065 ;
        RECT 104.705 219.765 105.590 219.935 ;
        RECT 103.550 219.085 104.060 219.175 ;
        RECT 102.100 218.275 102.325 218.405 ;
        RECT 102.495 218.335 103.020 218.555 ;
        RECT 103.190 218.915 104.060 219.085 ;
        RECT 101.735 217.685 101.985 218.145 ;
        RECT 102.155 218.135 102.325 218.275 ;
        RECT 103.190 218.135 103.360 218.915 ;
        RECT 103.890 218.845 104.060 218.915 ;
        RECT 103.570 218.665 103.770 218.695 ;
        RECT 104.230 218.665 104.400 219.735 ;
        RECT 104.570 218.845 104.760 219.565 ;
        RECT 103.570 218.365 104.400 218.665 ;
        RECT 104.930 218.635 105.250 219.595 ;
        RECT 102.155 217.965 102.490 218.135 ;
        RECT 102.685 217.965 103.360 218.135 ;
        RECT 103.680 217.685 104.050 218.185 ;
        RECT 104.230 218.135 104.400 218.365 ;
        RECT 104.785 218.305 105.250 218.635 ;
        RECT 105.420 218.925 105.590 219.765 ;
        RECT 105.770 219.735 106.085 220.235 ;
        RECT 106.315 219.505 106.655 220.065 ;
        RECT 105.760 219.130 106.655 219.505 ;
        RECT 106.825 219.225 106.995 220.235 ;
        RECT 106.465 218.925 106.655 219.130 ;
        RECT 107.165 219.175 107.495 220.020 ;
        RECT 107.785 219.175 108.115 220.020 ;
        RECT 108.285 219.225 108.455 220.235 ;
        RECT 108.625 219.505 108.965 220.065 ;
        RECT 109.195 219.735 109.510 220.235 ;
        RECT 109.690 219.765 110.575 219.935 ;
        RECT 107.165 219.095 107.555 219.175 ;
        RECT 107.340 219.045 107.555 219.095 ;
        RECT 105.420 218.595 106.295 218.925 ;
        RECT 106.465 218.595 107.215 218.925 ;
        RECT 105.420 218.135 105.590 218.595 ;
        RECT 106.465 218.425 106.665 218.595 ;
        RECT 107.385 218.465 107.555 219.045 ;
        RECT 107.330 218.425 107.555 218.465 ;
        RECT 104.230 217.965 104.635 218.135 ;
        RECT 104.805 217.965 105.590 218.135 ;
        RECT 105.865 217.685 106.075 218.215 ;
        RECT 106.335 217.900 106.665 218.425 ;
        RECT 107.175 218.340 107.555 218.425 ;
        RECT 107.725 219.095 108.115 219.175 ;
        RECT 108.625 219.130 109.520 219.505 ;
        RECT 107.725 219.045 107.940 219.095 ;
        RECT 107.725 218.465 107.895 219.045 ;
        RECT 108.625 218.925 108.815 219.130 ;
        RECT 109.690 218.925 109.860 219.765 ;
        RECT 110.800 219.735 111.050 220.065 ;
        RECT 108.065 218.595 108.815 218.925 ;
        RECT 108.985 218.595 109.860 218.925 ;
        RECT 107.725 218.425 107.950 218.465 ;
        RECT 108.615 218.425 108.815 218.595 ;
        RECT 107.725 218.340 108.105 218.425 ;
        RECT 106.835 217.685 107.005 218.295 ;
        RECT 107.175 217.905 107.505 218.340 ;
        RECT 107.775 217.905 108.105 218.340 ;
        RECT 108.275 217.685 108.445 218.295 ;
        RECT 108.615 217.900 108.945 218.425 ;
        RECT 109.205 217.685 109.415 218.215 ;
        RECT 109.690 218.135 109.860 218.595 ;
        RECT 110.030 218.635 110.350 219.595 ;
        RECT 110.520 218.845 110.710 219.565 ;
        RECT 110.880 218.665 111.050 219.735 ;
        RECT 111.220 219.435 111.390 220.235 ;
        RECT 111.560 219.790 112.665 219.960 ;
        RECT 111.560 219.175 111.730 219.790 ;
        RECT 112.875 219.640 113.125 220.065 ;
        RECT 113.295 219.775 113.560 220.235 ;
        RECT 111.900 219.255 112.430 219.620 ;
        RECT 112.875 219.510 113.180 219.640 ;
        RECT 111.220 219.085 111.730 219.175 ;
        RECT 111.220 218.915 112.090 219.085 ;
        RECT 111.220 218.845 111.390 218.915 ;
        RECT 111.510 218.665 111.710 218.695 ;
        RECT 110.030 218.305 110.495 218.635 ;
        RECT 110.880 218.365 111.710 218.665 ;
        RECT 110.880 218.135 111.050 218.365 ;
        RECT 109.690 217.965 110.475 218.135 ;
        RECT 110.645 217.965 111.050 218.135 ;
        RECT 111.230 217.685 111.600 218.185 ;
        RECT 111.920 218.135 112.090 218.915 ;
        RECT 112.260 218.555 112.430 219.255 ;
        RECT 112.600 218.725 112.840 219.320 ;
        RECT 112.260 218.335 112.785 218.555 ;
        RECT 113.010 218.405 113.180 219.510 ;
        RECT 112.955 218.275 113.180 218.405 ;
        RECT 113.350 218.315 113.630 219.265 ;
        RECT 112.955 218.135 113.125 218.275 ;
        RECT 111.920 217.965 112.595 218.135 ;
        RECT 112.790 217.965 113.125 218.135 ;
        RECT 113.295 217.685 113.545 218.145 ;
        RECT 113.800 217.945 113.985 220.065 ;
        RECT 114.155 219.735 114.485 220.235 ;
        RECT 114.655 219.565 114.825 220.065 ;
        RECT 114.160 219.395 114.825 219.565 ;
        RECT 115.105 219.645 115.345 220.035 ;
        RECT 115.515 219.825 115.865 220.235 ;
        RECT 115.105 219.445 115.855 219.645 ;
        RECT 114.160 218.405 114.390 219.395 ;
        RECT 114.560 218.575 114.910 219.225 ;
        RECT 114.160 218.235 114.825 218.405 ;
        RECT 114.155 217.685 114.485 218.065 ;
        RECT 114.655 217.945 114.825 218.235 ;
        RECT 115.105 217.925 115.335 219.265 ;
        RECT 115.515 218.765 115.855 219.445 ;
        RECT 116.035 218.945 116.365 220.055 ;
        RECT 116.535 219.585 116.715 220.055 ;
        RECT 116.885 219.755 117.215 220.235 ;
        RECT 117.390 219.585 117.560 220.055 ;
        RECT 116.535 219.385 117.560 219.585 ;
        RECT 115.515 217.865 115.745 218.765 ;
        RECT 116.035 218.645 116.580 218.945 ;
        RECT 115.945 217.685 116.190 218.465 ;
        RECT 116.360 218.415 116.580 218.645 ;
        RECT 116.750 218.595 117.175 219.215 ;
        RECT 117.370 218.595 117.630 219.215 ;
        RECT 117.825 219.095 118.110 220.235 ;
        RECT 117.840 218.415 118.100 218.925 ;
        RECT 116.360 218.225 118.100 218.415 ;
        RECT 116.360 217.865 116.790 218.225 ;
        RECT 117.370 217.685 118.100 218.055 ;
        RECT 118.300 217.865 118.580 220.055 ;
        RECT 118.765 219.070 119.055 220.235 ;
        RECT 119.285 219.095 119.495 220.235 ;
        RECT 119.665 219.085 119.995 220.065 ;
        RECT 120.165 219.095 120.395 220.235 ;
        RECT 121.615 219.565 121.785 220.065 ;
        RECT 121.955 219.735 122.285 220.235 ;
        RECT 121.615 219.395 122.280 219.565 ;
        RECT 118.765 217.685 119.055 218.410 ;
        RECT 119.285 217.685 119.495 218.505 ;
        RECT 119.665 218.485 119.915 219.085 ;
        RECT 120.085 218.675 120.415 218.925 ;
        RECT 121.530 218.575 121.880 219.225 ;
        RECT 119.665 217.855 119.995 218.485 ;
        RECT 120.165 217.685 120.395 218.505 ;
        RECT 122.050 218.405 122.280 219.395 ;
        RECT 121.615 218.235 122.280 218.405 ;
        RECT 121.615 217.945 121.785 218.235 ;
        RECT 121.955 217.685 122.285 218.065 ;
        RECT 122.455 217.945 122.640 220.065 ;
        RECT 122.880 219.775 123.145 220.235 ;
        RECT 123.315 219.640 123.565 220.065 ;
        RECT 123.775 219.790 124.880 219.960 ;
        RECT 123.260 219.510 123.565 219.640 ;
        RECT 122.810 218.315 123.090 219.265 ;
        RECT 123.260 218.405 123.430 219.510 ;
        RECT 123.600 218.725 123.840 219.320 ;
        RECT 124.010 219.255 124.540 219.620 ;
        RECT 124.010 218.555 124.180 219.255 ;
        RECT 124.710 219.175 124.880 219.790 ;
        RECT 125.050 219.435 125.220 220.235 ;
        RECT 125.390 219.735 125.640 220.065 ;
        RECT 125.865 219.765 126.750 219.935 ;
        RECT 124.710 219.085 125.220 219.175 ;
        RECT 123.260 218.275 123.485 218.405 ;
        RECT 123.655 218.335 124.180 218.555 ;
        RECT 124.350 218.915 125.220 219.085 ;
        RECT 122.895 217.685 123.145 218.145 ;
        RECT 123.315 218.135 123.485 218.275 ;
        RECT 124.350 218.135 124.520 218.915 ;
        RECT 125.050 218.845 125.220 218.915 ;
        RECT 124.730 218.665 124.930 218.695 ;
        RECT 125.390 218.665 125.560 219.735 ;
        RECT 125.730 218.845 125.920 219.565 ;
        RECT 124.730 218.365 125.560 218.665 ;
        RECT 126.090 218.635 126.410 219.595 ;
        RECT 123.315 217.965 123.650 218.135 ;
        RECT 123.845 217.965 124.520 218.135 ;
        RECT 124.840 217.685 125.210 218.185 ;
        RECT 125.390 218.135 125.560 218.365 ;
        RECT 125.945 218.305 126.410 218.635 ;
        RECT 126.580 218.925 126.750 219.765 ;
        RECT 126.930 219.735 127.245 220.235 ;
        RECT 127.475 219.505 127.815 220.065 ;
        RECT 126.920 219.130 127.815 219.505 ;
        RECT 127.985 219.225 128.155 220.235 ;
        RECT 127.625 218.925 127.815 219.130 ;
        RECT 128.325 219.175 128.655 220.020 ;
        RECT 128.325 219.095 128.715 219.175 ;
        RECT 128.885 219.145 132.395 220.235 ;
        RECT 133.115 219.565 133.285 220.065 ;
        RECT 133.455 219.735 133.785 220.235 ;
        RECT 133.115 219.395 133.780 219.565 ;
        RECT 128.500 219.045 128.715 219.095 ;
        RECT 126.580 218.595 127.455 218.925 ;
        RECT 127.625 218.595 128.375 218.925 ;
        RECT 126.580 218.135 126.750 218.595 ;
        RECT 127.625 218.425 127.825 218.595 ;
        RECT 128.545 218.465 128.715 219.045 ;
        RECT 128.490 218.445 128.715 218.465 ;
        RECT 128.485 218.425 128.715 218.445 ;
        RECT 125.390 217.965 125.795 218.135 ;
        RECT 125.965 217.965 126.750 218.135 ;
        RECT 127.025 217.685 127.235 218.215 ;
        RECT 127.495 217.900 127.825 218.425 ;
        RECT 128.335 218.340 128.715 218.425 ;
        RECT 128.885 218.455 130.535 218.975 ;
        RECT 130.705 218.625 132.395 219.145 ;
        RECT 133.030 218.575 133.380 219.225 ;
        RECT 127.995 217.685 128.165 218.295 ;
        RECT 128.335 217.905 128.665 218.340 ;
        RECT 128.885 217.685 132.395 218.455 ;
        RECT 133.550 218.405 133.780 219.395 ;
        RECT 133.115 218.235 133.780 218.405 ;
        RECT 133.115 217.945 133.285 218.235 ;
        RECT 133.455 217.685 133.785 218.065 ;
        RECT 133.955 217.945 134.140 220.065 ;
        RECT 134.380 219.775 134.645 220.235 ;
        RECT 134.815 219.640 135.065 220.065 ;
        RECT 135.275 219.790 136.380 219.960 ;
        RECT 134.760 219.510 135.065 219.640 ;
        RECT 134.310 218.315 134.590 219.265 ;
        RECT 134.760 218.405 134.930 219.510 ;
        RECT 135.100 218.725 135.340 219.320 ;
        RECT 135.510 219.255 136.040 219.620 ;
        RECT 135.510 218.555 135.680 219.255 ;
        RECT 136.210 219.175 136.380 219.790 ;
        RECT 136.550 219.435 136.720 220.235 ;
        RECT 136.890 219.735 137.140 220.065 ;
        RECT 137.365 219.765 138.250 219.935 ;
        RECT 136.210 219.085 136.720 219.175 ;
        RECT 134.760 218.275 134.985 218.405 ;
        RECT 135.155 218.335 135.680 218.555 ;
        RECT 135.850 218.915 136.720 219.085 ;
        RECT 134.395 217.685 134.645 218.145 ;
        RECT 134.815 218.135 134.985 218.275 ;
        RECT 135.850 218.135 136.020 218.915 ;
        RECT 136.550 218.845 136.720 218.915 ;
        RECT 136.230 218.665 136.430 218.695 ;
        RECT 136.890 218.665 137.060 219.735 ;
        RECT 137.230 218.845 137.420 219.565 ;
        RECT 136.230 218.365 137.060 218.665 ;
        RECT 137.590 218.635 137.910 219.595 ;
        RECT 134.815 217.965 135.150 218.135 ;
        RECT 135.345 217.965 136.020 218.135 ;
        RECT 136.340 217.685 136.710 218.185 ;
        RECT 136.890 218.135 137.060 218.365 ;
        RECT 137.445 218.305 137.910 218.635 ;
        RECT 138.080 218.925 138.250 219.765 ;
        RECT 138.430 219.735 138.745 220.235 ;
        RECT 138.975 219.505 139.315 220.065 ;
        RECT 138.420 219.130 139.315 219.505 ;
        RECT 139.485 219.225 139.655 220.235 ;
        RECT 139.125 218.925 139.315 219.130 ;
        RECT 139.825 219.175 140.155 220.020 ;
        RECT 140.385 219.475 140.900 219.885 ;
        RECT 141.135 219.475 141.305 220.235 ;
        RECT 141.475 219.895 143.505 220.065 ;
        RECT 139.825 219.095 140.215 219.175 ;
        RECT 140.000 219.045 140.215 219.095 ;
        RECT 138.080 218.595 138.955 218.925 ;
        RECT 139.125 218.595 139.875 218.925 ;
        RECT 138.080 218.135 138.250 218.595 ;
        RECT 139.125 218.425 139.325 218.595 ;
        RECT 140.045 218.465 140.215 219.045 ;
        RECT 140.385 218.665 140.725 219.475 ;
        RECT 141.475 219.230 141.645 219.895 ;
        RECT 142.040 219.555 143.165 219.725 ;
        RECT 140.895 219.040 141.645 219.230 ;
        RECT 141.815 219.215 142.825 219.385 ;
        RECT 140.905 218.955 141.075 219.040 ;
        RECT 140.385 218.495 141.615 218.665 ;
        RECT 139.990 218.445 140.215 218.465 ;
        RECT 139.985 218.425 140.215 218.445 ;
        RECT 136.890 217.965 137.295 218.135 ;
        RECT 137.465 217.965 138.250 218.135 ;
        RECT 138.525 217.685 138.735 218.215 ;
        RECT 138.995 217.900 139.325 218.425 ;
        RECT 139.835 218.340 140.215 218.425 ;
        RECT 139.495 217.685 139.665 218.295 ;
        RECT 139.835 217.905 140.165 218.340 ;
        RECT 140.660 217.890 140.905 218.495 ;
        RECT 141.125 217.685 141.635 218.220 ;
        RECT 141.815 217.855 142.005 219.215 ;
        RECT 142.175 218.445 142.450 219.015 ;
        RECT 142.175 218.275 142.455 218.445 ;
        RECT 142.655 218.415 142.825 219.215 ;
        RECT 142.995 218.425 143.165 219.555 ;
        RECT 143.335 218.925 143.505 219.895 ;
        RECT 143.675 219.095 143.845 220.235 ;
        RECT 144.015 219.095 144.350 220.065 ;
        RECT 143.335 218.595 143.530 218.925 ;
        RECT 143.755 218.595 144.010 218.925 ;
        RECT 143.755 218.425 143.925 218.595 ;
        RECT 144.180 218.445 144.350 219.095 ;
        RECT 144.525 219.070 144.815 220.235 ;
        RECT 145.075 219.565 145.245 220.065 ;
        RECT 145.415 219.735 145.745 220.235 ;
        RECT 145.075 219.395 145.740 219.565 ;
        RECT 144.990 218.575 145.340 219.225 ;
        RECT 144.125 218.425 144.350 218.445 ;
        RECT 142.175 217.855 142.450 218.275 ;
        RECT 142.995 218.255 143.925 218.425 ;
        RECT 142.995 218.220 143.170 218.255 ;
        RECT 142.640 217.855 143.170 218.220 ;
        RECT 143.595 217.685 143.925 218.085 ;
        RECT 144.095 217.855 144.350 218.425 ;
        RECT 144.525 217.685 144.815 218.410 ;
        RECT 145.510 218.405 145.740 219.395 ;
        RECT 145.075 218.235 145.740 218.405 ;
        RECT 145.075 217.945 145.245 218.235 ;
        RECT 145.415 217.685 145.745 218.065 ;
        RECT 145.915 217.945 146.100 220.065 ;
        RECT 146.340 219.775 146.605 220.235 ;
        RECT 146.775 219.640 147.025 220.065 ;
        RECT 147.235 219.790 148.340 219.960 ;
        RECT 146.720 219.510 147.025 219.640 ;
        RECT 146.270 218.315 146.550 219.265 ;
        RECT 146.720 218.405 146.890 219.510 ;
        RECT 147.060 218.725 147.300 219.320 ;
        RECT 147.470 219.255 148.000 219.620 ;
        RECT 147.470 218.555 147.640 219.255 ;
        RECT 148.170 219.175 148.340 219.790 ;
        RECT 148.510 219.435 148.680 220.235 ;
        RECT 148.850 219.735 149.100 220.065 ;
        RECT 149.325 219.765 150.210 219.935 ;
        RECT 148.170 219.085 148.680 219.175 ;
        RECT 146.720 218.275 146.945 218.405 ;
        RECT 147.115 218.335 147.640 218.555 ;
        RECT 147.810 218.915 148.680 219.085 ;
        RECT 146.355 217.685 146.605 218.145 ;
        RECT 146.775 218.135 146.945 218.275 ;
        RECT 147.810 218.135 147.980 218.915 ;
        RECT 148.510 218.845 148.680 218.915 ;
        RECT 148.190 218.665 148.390 218.695 ;
        RECT 148.850 218.665 149.020 219.735 ;
        RECT 149.190 218.845 149.380 219.565 ;
        RECT 148.190 218.365 149.020 218.665 ;
        RECT 149.550 218.635 149.870 219.595 ;
        RECT 146.775 217.965 147.110 218.135 ;
        RECT 147.305 217.965 147.980 218.135 ;
        RECT 148.300 217.685 148.670 218.185 ;
        RECT 148.850 218.135 149.020 218.365 ;
        RECT 149.405 218.305 149.870 218.635 ;
        RECT 150.040 218.925 150.210 219.765 ;
        RECT 150.390 219.735 150.705 220.235 ;
        RECT 150.935 219.505 151.275 220.065 ;
        RECT 150.380 219.130 151.275 219.505 ;
        RECT 151.445 219.225 151.615 220.235 ;
        RECT 151.085 218.925 151.275 219.130 ;
        RECT 151.785 219.175 152.115 220.020 ;
        RECT 151.785 219.095 152.175 219.175 ;
        RECT 151.960 219.045 152.175 219.095 ;
        RECT 150.040 218.595 150.915 218.925 ;
        RECT 151.085 218.595 151.835 218.925 ;
        RECT 150.040 218.135 150.210 218.595 ;
        RECT 151.085 218.425 151.285 218.595 ;
        RECT 152.005 218.465 152.175 219.045 ;
        RECT 151.950 218.425 152.175 218.465 ;
        RECT 148.850 217.965 149.255 218.135 ;
        RECT 149.425 217.965 150.210 218.135 ;
        RECT 150.485 217.685 150.695 218.215 ;
        RECT 150.955 217.900 151.285 218.425 ;
        RECT 151.795 218.340 152.175 218.425 ;
        RECT 152.805 219.095 153.190 220.065 ;
        RECT 153.360 219.775 153.685 220.235 ;
        RECT 154.205 219.605 154.485 220.065 ;
        RECT 153.360 219.385 154.485 219.605 ;
        RECT 152.805 218.425 153.085 219.095 ;
        RECT 153.360 218.925 153.810 219.385 ;
        RECT 154.675 219.215 155.075 220.065 ;
        RECT 155.475 219.775 155.745 220.235 ;
        RECT 155.915 219.605 156.200 220.065 ;
        RECT 153.255 218.595 153.810 218.925 ;
        RECT 153.980 218.655 155.075 219.215 ;
        RECT 153.360 218.485 153.810 218.595 ;
        RECT 151.455 217.685 151.625 218.295 ;
        RECT 151.795 217.905 152.125 218.340 ;
        RECT 152.805 217.855 153.190 218.425 ;
        RECT 153.360 218.315 154.485 218.485 ;
        RECT 153.360 217.685 153.685 218.145 ;
        RECT 154.205 217.855 154.485 218.315 ;
        RECT 154.675 217.855 155.075 218.655 ;
        RECT 155.245 219.385 156.200 219.605 ;
        RECT 155.245 218.485 155.455 219.385 ;
        RECT 155.625 218.655 156.315 219.215 ;
        RECT 156.945 219.145 158.155 220.235 ;
        RECT 156.945 218.605 157.465 219.145 ;
        RECT 155.245 218.315 156.200 218.485 ;
        RECT 157.635 218.435 158.155 218.975 ;
        RECT 155.475 217.685 155.745 218.145 ;
        RECT 155.915 217.855 156.200 218.315 ;
        RECT 156.945 217.685 158.155 218.435 ;
        RECT 2.760 217.515 158.240 217.685 ;
        RECT 2.845 216.765 4.055 217.515 ;
        RECT 4.225 216.970 9.570 217.515 ;
        RECT 9.745 216.970 15.090 217.515 ;
        RECT 15.265 216.970 20.610 217.515 ;
        RECT 20.785 216.970 26.130 217.515 ;
        RECT 2.845 216.225 3.365 216.765 ;
        RECT 3.535 216.055 4.055 216.595 ;
        RECT 5.810 216.140 6.150 216.970 ;
        RECT 2.845 214.965 4.055 216.055 ;
        RECT 7.630 215.400 7.980 216.650 ;
        RECT 11.330 216.140 11.670 216.970 ;
        RECT 13.150 215.400 13.500 216.650 ;
        RECT 16.850 216.140 17.190 216.970 ;
        RECT 18.670 215.400 19.020 216.650 ;
        RECT 22.370 216.140 22.710 216.970 ;
        RECT 26.305 216.745 27.975 217.515 ;
        RECT 28.605 216.790 28.895 217.515 ;
        RECT 29.065 216.970 34.410 217.515 ;
        RECT 34.585 216.970 39.930 217.515 ;
        RECT 40.105 216.970 45.450 217.515 ;
        RECT 45.625 216.970 50.970 217.515 ;
        RECT 24.190 215.400 24.540 216.650 ;
        RECT 26.305 216.225 27.055 216.745 ;
        RECT 27.225 216.055 27.975 216.575 ;
        RECT 30.650 216.140 30.990 216.970 ;
        RECT 4.225 214.965 9.570 215.400 ;
        RECT 9.745 214.965 15.090 215.400 ;
        RECT 15.265 214.965 20.610 215.400 ;
        RECT 20.785 214.965 26.130 215.400 ;
        RECT 26.305 214.965 27.975 216.055 ;
        RECT 28.605 214.965 28.895 216.130 ;
        RECT 32.470 215.400 32.820 216.650 ;
        RECT 36.170 216.140 36.510 216.970 ;
        RECT 37.990 215.400 38.340 216.650 ;
        RECT 41.690 216.140 42.030 216.970 ;
        RECT 43.510 215.400 43.860 216.650 ;
        RECT 47.210 216.140 47.550 216.970 ;
        RECT 51.145 216.745 53.735 217.515 ;
        RECT 54.365 216.790 54.655 217.515 ;
        RECT 54.825 216.745 56.495 217.515 ;
        RECT 56.755 217.035 57.055 217.515 ;
        RECT 57.225 216.865 57.485 217.320 ;
        RECT 57.655 217.035 57.915 217.515 ;
        RECT 58.095 216.865 58.355 217.320 ;
        RECT 58.525 217.035 58.775 217.515 ;
        RECT 58.955 216.865 59.215 217.320 ;
        RECT 59.385 217.035 59.635 217.515 ;
        RECT 59.815 216.865 60.075 217.320 ;
        RECT 60.245 217.035 60.490 217.515 ;
        RECT 60.660 216.865 60.935 217.320 ;
        RECT 61.105 217.035 61.350 217.515 ;
        RECT 61.520 216.865 61.780 217.320 ;
        RECT 61.950 217.035 62.210 217.515 ;
        RECT 62.380 216.865 62.640 217.320 ;
        RECT 62.810 217.035 63.070 217.515 ;
        RECT 63.240 216.865 63.500 217.320 ;
        RECT 63.670 216.955 63.930 217.515 ;
        RECT 49.030 215.400 49.380 216.650 ;
        RECT 51.145 216.225 52.355 216.745 ;
        RECT 52.525 216.055 53.735 216.575 ;
        RECT 54.825 216.225 55.575 216.745 ;
        RECT 56.755 216.695 63.500 216.865 ;
        RECT 29.065 214.965 34.410 215.400 ;
        RECT 34.585 214.965 39.930 215.400 ;
        RECT 40.105 214.965 45.450 215.400 ;
        RECT 45.625 214.965 50.970 215.400 ;
        RECT 51.145 214.965 53.735 216.055 ;
        RECT 54.365 214.965 54.655 216.130 ;
        RECT 55.745 216.055 56.495 216.575 ;
        RECT 56.755 216.105 57.920 216.695 ;
        RECT 64.100 216.525 64.350 217.335 ;
        RECT 64.530 216.990 64.790 217.515 ;
        RECT 64.960 216.525 65.210 217.335 ;
        RECT 65.390 217.005 65.695 217.515 ;
        RECT 65.925 217.055 66.170 217.515 ;
        RECT 58.090 216.275 65.210 216.525 ;
        RECT 65.380 216.275 65.695 216.835 ;
        RECT 65.865 216.275 66.180 216.885 ;
        RECT 66.350 216.525 66.600 217.335 ;
        RECT 66.770 216.990 67.030 217.515 ;
        RECT 67.200 216.865 67.460 217.320 ;
        RECT 67.630 217.035 67.890 217.515 ;
        RECT 68.060 216.865 68.320 217.320 ;
        RECT 68.490 217.035 68.750 217.515 ;
        RECT 68.920 216.865 69.180 217.320 ;
        RECT 69.350 217.035 69.610 217.515 ;
        RECT 69.780 216.865 70.040 217.320 ;
        RECT 70.210 217.035 70.510 217.515 ;
        RECT 70.930 217.260 71.265 217.305 ;
        RECT 67.200 216.695 70.510 216.865 ;
        RECT 66.350 216.275 69.370 216.525 ;
        RECT 56.755 216.065 63.500 216.105 ;
        RECT 54.825 214.965 56.495 216.055 ;
        RECT 56.725 215.895 63.500 216.065 ;
        RECT 56.755 215.880 63.500 215.895 ;
        RECT 56.755 214.965 57.025 215.710 ;
        RECT 57.195 215.140 57.485 215.880 ;
        RECT 58.095 215.865 63.500 215.880 ;
        RECT 57.655 214.970 57.910 215.695 ;
        RECT 58.095 215.140 58.355 215.865 ;
        RECT 58.525 214.970 58.770 215.695 ;
        RECT 58.955 215.140 59.215 215.865 ;
        RECT 59.385 214.970 59.630 215.695 ;
        RECT 59.815 215.140 60.075 215.865 ;
        RECT 60.245 214.970 60.490 215.695 ;
        RECT 60.660 215.140 60.920 215.865 ;
        RECT 61.090 214.970 61.350 215.695 ;
        RECT 61.520 215.140 61.780 215.865 ;
        RECT 61.950 214.970 62.210 215.695 ;
        RECT 62.380 215.140 62.640 215.865 ;
        RECT 62.810 214.970 63.070 215.695 ;
        RECT 63.240 215.140 63.500 215.865 ;
        RECT 63.670 214.970 63.930 215.765 ;
        RECT 64.100 215.140 64.350 216.275 ;
        RECT 57.655 214.965 63.930 214.970 ;
        RECT 64.530 214.965 64.790 215.775 ;
        RECT 64.965 215.135 65.210 216.275 ;
        RECT 65.465 216.235 65.635 216.275 ;
        RECT 65.390 214.965 65.685 215.775 ;
        RECT 65.875 214.965 66.170 216.075 ;
        RECT 66.350 215.140 66.600 216.275 ;
        RECT 69.540 216.105 70.510 216.695 ;
        RECT 66.770 214.965 67.030 216.075 ;
        RECT 67.200 215.865 70.510 216.105 ;
        RECT 70.925 216.795 71.265 217.260 ;
        RECT 71.435 217.135 71.765 217.515 ;
        RECT 72.225 217.085 72.495 217.180 ;
        RECT 70.925 216.105 71.095 216.795 ;
        RECT 71.265 216.275 71.525 216.605 ;
        RECT 67.200 215.140 67.460 215.865 ;
        RECT 67.630 214.965 67.890 215.695 ;
        RECT 68.060 215.140 68.320 215.865 ;
        RECT 68.490 214.965 68.750 215.695 ;
        RECT 68.920 215.140 69.180 215.865 ;
        RECT 69.350 214.965 69.610 215.695 ;
        RECT 69.780 215.140 70.040 215.865 ;
        RECT 70.210 214.965 70.505 215.695 ;
        RECT 70.925 215.135 71.185 216.105 ;
        RECT 71.355 215.725 71.525 216.275 ;
        RECT 71.695 215.905 72.035 216.935 ;
        RECT 72.225 216.915 72.535 217.085 ;
        RECT 72.225 215.905 72.495 216.915 ;
        RECT 72.720 215.905 73.000 217.180 ;
        RECT 73.200 217.015 73.430 217.345 ;
        RECT 73.675 217.135 74.005 217.515 ;
        RECT 72.825 215.895 72.995 215.905 ;
        RECT 73.200 215.725 73.370 217.015 ;
        RECT 74.175 216.945 74.350 217.345 ;
        RECT 75.085 217.045 75.380 217.515 ;
        RECT 73.720 216.775 74.350 216.945 ;
        RECT 75.550 216.875 75.810 217.320 ;
        RECT 75.980 217.045 76.240 217.515 ;
        RECT 76.410 216.875 76.665 217.320 ;
        RECT 76.835 217.045 77.135 217.515 ;
        RECT 73.720 216.605 73.890 216.775 ;
        RECT 74.625 216.705 77.655 216.875 ;
        RECT 73.540 216.275 73.890 216.605 ;
        RECT 71.355 215.555 73.370 215.725 ;
        RECT 73.720 215.755 73.890 216.275 ;
        RECT 74.070 215.925 74.435 216.605 ;
        RECT 74.625 216.140 74.795 216.705 ;
        RECT 74.965 216.310 77.180 216.535 ;
        RECT 77.355 216.140 77.655 216.705 ;
        RECT 78.785 216.695 79.015 217.515 ;
        RECT 79.185 216.715 79.515 217.345 ;
        RECT 78.765 216.275 79.095 216.525 ;
        RECT 74.625 215.970 77.655 216.140 ;
        RECT 79.265 216.115 79.515 216.715 ;
        RECT 79.685 216.695 79.895 217.515 ;
        RECT 80.125 216.790 80.415 217.515 ;
        RECT 80.675 216.965 80.845 217.255 ;
        RECT 81.015 217.135 81.345 217.515 ;
        RECT 80.675 216.795 81.340 216.965 ;
        RECT 73.720 215.585 74.350 215.755 ;
        RECT 71.380 214.965 71.710 215.375 ;
        RECT 71.910 215.135 72.080 215.555 ;
        RECT 72.295 214.965 72.965 215.375 ;
        RECT 73.200 215.135 73.370 215.555 ;
        RECT 73.675 214.965 74.005 215.405 ;
        RECT 74.175 215.135 74.350 215.585 ;
        RECT 74.605 214.965 74.950 215.800 ;
        RECT 75.125 215.165 75.380 215.970 ;
        RECT 75.550 214.965 75.810 215.800 ;
        RECT 75.985 215.165 76.240 215.970 ;
        RECT 76.410 214.965 76.670 215.800 ;
        RECT 76.840 215.165 77.100 215.970 ;
        RECT 77.270 214.965 77.655 215.800 ;
        RECT 78.785 214.965 79.015 216.105 ;
        RECT 79.185 215.135 79.515 216.115 ;
        RECT 79.685 214.965 79.895 216.105 ;
        RECT 80.125 214.965 80.415 216.130 ;
        RECT 80.590 215.975 80.940 216.625 ;
        RECT 81.110 215.805 81.340 216.795 ;
        RECT 80.675 215.635 81.340 215.805 ;
        RECT 80.675 215.135 80.845 215.635 ;
        RECT 81.015 214.965 81.345 215.465 ;
        RECT 81.515 215.135 81.700 217.255 ;
        RECT 81.955 217.055 82.205 217.515 ;
        RECT 82.375 217.065 82.710 217.235 ;
        RECT 82.905 217.065 83.580 217.235 ;
        RECT 82.375 216.925 82.545 217.065 ;
        RECT 81.870 215.935 82.150 216.885 ;
        RECT 82.320 216.795 82.545 216.925 ;
        RECT 82.320 215.690 82.490 216.795 ;
        RECT 82.715 216.645 83.240 216.865 ;
        RECT 82.660 215.880 82.900 216.475 ;
        RECT 83.070 215.945 83.240 216.645 ;
        RECT 83.410 216.285 83.580 217.065 ;
        RECT 83.900 217.015 84.270 217.515 ;
        RECT 84.450 217.065 84.855 217.235 ;
        RECT 85.025 217.065 85.810 217.235 ;
        RECT 84.450 216.835 84.620 217.065 ;
        RECT 83.790 216.535 84.620 216.835 ;
        RECT 85.005 216.565 85.470 216.895 ;
        RECT 83.790 216.505 83.990 216.535 ;
        RECT 84.110 216.285 84.280 216.355 ;
        RECT 83.410 216.115 84.280 216.285 ;
        RECT 83.770 216.025 84.280 216.115 ;
        RECT 82.320 215.560 82.625 215.690 ;
        RECT 83.070 215.580 83.600 215.945 ;
        RECT 81.940 214.965 82.205 215.425 ;
        RECT 82.375 215.135 82.625 215.560 ;
        RECT 83.770 215.410 83.940 216.025 ;
        RECT 82.835 215.240 83.940 215.410 ;
        RECT 84.110 214.965 84.280 215.765 ;
        RECT 84.450 215.465 84.620 216.535 ;
        RECT 84.790 215.635 84.980 216.355 ;
        RECT 85.150 215.605 85.470 216.565 ;
        RECT 85.640 216.605 85.810 217.065 ;
        RECT 86.085 216.985 86.295 217.515 ;
        RECT 86.555 216.775 86.885 217.300 ;
        RECT 87.055 216.905 87.225 217.515 ;
        RECT 87.395 216.860 87.725 217.295 ;
        RECT 88.115 217.000 88.285 217.515 ;
        RECT 88.455 216.860 88.785 217.295 ;
        RECT 88.955 216.905 89.125 217.515 ;
        RECT 87.395 216.775 87.775 216.860 ;
        RECT 86.685 216.605 86.885 216.775 ;
        RECT 87.550 216.735 87.775 216.775 ;
        RECT 85.640 216.275 86.515 216.605 ;
        RECT 86.685 216.275 87.435 216.605 ;
        RECT 84.450 215.135 84.700 215.465 ;
        RECT 85.640 215.435 85.810 216.275 ;
        RECT 86.685 216.070 86.875 216.275 ;
        RECT 87.605 216.155 87.775 216.735 ;
        RECT 87.560 216.105 87.775 216.155 ;
        RECT 85.980 215.695 86.875 216.070 ;
        RECT 87.385 216.025 87.775 216.105 ;
        RECT 88.405 216.775 88.785 216.860 ;
        RECT 89.295 216.775 89.625 217.300 ;
        RECT 89.885 216.985 90.095 217.515 ;
        RECT 90.370 217.065 91.155 217.235 ;
        RECT 91.325 217.065 91.730 217.235 ;
        RECT 88.405 216.735 88.630 216.775 ;
        RECT 88.405 216.155 88.575 216.735 ;
        RECT 89.295 216.605 89.495 216.775 ;
        RECT 90.370 216.605 90.540 217.065 ;
        RECT 88.745 216.275 89.495 216.605 ;
        RECT 89.665 216.275 90.540 216.605 ;
        RECT 88.405 216.105 88.620 216.155 ;
        RECT 88.405 216.025 88.795 216.105 ;
        RECT 84.925 215.265 85.810 215.435 ;
        RECT 85.990 214.965 86.305 215.465 ;
        RECT 86.535 215.135 86.875 215.695 ;
        RECT 87.045 214.965 87.215 215.975 ;
        RECT 87.385 215.180 87.715 216.025 ;
        RECT 88.125 214.965 88.295 215.880 ;
        RECT 88.465 215.180 88.795 216.025 ;
        RECT 89.305 216.070 89.495 216.275 ;
        RECT 88.965 214.965 89.135 215.975 ;
        RECT 89.305 215.695 90.200 216.070 ;
        RECT 89.305 215.135 89.645 215.695 ;
        RECT 89.875 214.965 90.190 215.465 ;
        RECT 90.370 215.435 90.540 216.275 ;
        RECT 90.710 216.565 91.175 216.895 ;
        RECT 91.560 216.835 91.730 217.065 ;
        RECT 91.910 217.015 92.280 217.515 ;
        RECT 92.600 217.065 93.275 217.235 ;
        RECT 93.470 217.065 93.805 217.235 ;
        RECT 90.710 215.605 91.030 216.565 ;
        RECT 91.560 216.535 92.390 216.835 ;
        RECT 91.200 215.635 91.390 216.355 ;
        RECT 91.560 215.465 91.730 216.535 ;
        RECT 92.190 216.505 92.390 216.535 ;
        RECT 91.900 216.285 92.070 216.355 ;
        RECT 92.600 216.285 92.770 217.065 ;
        RECT 93.635 216.925 93.805 217.065 ;
        RECT 93.975 217.055 94.225 217.515 ;
        RECT 91.900 216.115 92.770 216.285 ;
        RECT 92.940 216.645 93.465 216.865 ;
        RECT 93.635 216.795 93.860 216.925 ;
        RECT 91.900 216.025 92.410 216.115 ;
        RECT 90.370 215.265 91.255 215.435 ;
        RECT 91.480 215.135 91.730 215.465 ;
        RECT 91.900 214.965 92.070 215.765 ;
        RECT 92.240 215.410 92.410 216.025 ;
        RECT 92.940 215.945 93.110 216.645 ;
        RECT 92.580 215.580 93.110 215.945 ;
        RECT 93.280 215.880 93.520 216.475 ;
        RECT 93.690 215.690 93.860 216.795 ;
        RECT 94.030 215.935 94.310 216.885 ;
        RECT 93.555 215.560 93.860 215.690 ;
        RECT 92.240 215.240 93.345 215.410 ;
        RECT 93.555 215.135 93.805 215.560 ;
        RECT 93.975 214.965 94.240 215.425 ;
        RECT 94.480 215.135 94.665 217.255 ;
        RECT 94.835 217.135 95.165 217.515 ;
        RECT 95.335 216.965 95.505 217.255 ;
        RECT 94.840 216.795 95.505 216.965 ;
        RECT 96.690 216.965 96.945 217.255 ;
        RECT 97.115 217.135 97.445 217.515 ;
        RECT 96.690 216.795 97.440 216.965 ;
        RECT 94.840 215.805 95.070 216.795 ;
        RECT 95.240 215.975 95.590 216.625 ;
        RECT 96.690 215.975 97.040 216.625 ;
        RECT 97.210 215.805 97.440 216.795 ;
        RECT 94.840 215.635 95.505 215.805 ;
        RECT 94.835 214.965 95.165 215.465 ;
        RECT 95.335 215.135 95.505 215.635 ;
        RECT 96.690 215.635 97.440 215.805 ;
        RECT 96.690 215.135 96.945 215.635 ;
        RECT 97.115 214.965 97.445 215.465 ;
        RECT 97.615 215.135 97.785 217.255 ;
        RECT 98.145 217.155 98.475 217.515 ;
        RECT 98.645 217.125 99.140 217.295 ;
        RECT 99.345 217.125 100.200 217.295 ;
        RECT 98.015 215.935 98.475 216.985 ;
        RECT 97.955 215.150 98.280 215.935 ;
        RECT 98.645 215.765 98.815 217.125 ;
        RECT 98.985 216.215 99.335 216.835 ;
        RECT 99.505 216.615 99.860 216.835 ;
        RECT 99.505 216.025 99.675 216.615 ;
        RECT 100.030 216.415 100.200 217.125 ;
        RECT 101.075 217.055 101.405 217.515 ;
        RECT 101.615 217.155 101.965 217.325 ;
        RECT 100.405 216.585 101.195 216.835 ;
        RECT 101.615 216.765 101.875 217.155 ;
        RECT 102.185 217.065 103.135 217.345 ;
        RECT 103.305 217.075 103.495 217.515 ;
        RECT 103.665 217.135 104.735 217.305 ;
        RECT 101.365 216.415 101.535 216.595 ;
        RECT 98.645 215.595 99.040 215.765 ;
        RECT 99.210 215.635 99.675 216.025 ;
        RECT 99.845 216.245 101.535 216.415 ;
        RECT 98.870 215.465 99.040 215.595 ;
        RECT 99.845 215.465 100.015 216.245 ;
        RECT 101.705 216.075 101.875 216.765 ;
        RECT 100.375 215.905 101.875 216.075 ;
        RECT 102.065 216.105 102.275 216.895 ;
        RECT 102.445 216.275 102.795 216.895 ;
        RECT 102.965 216.285 103.135 217.065 ;
        RECT 103.665 216.905 103.835 217.135 ;
        RECT 103.305 216.735 103.835 216.905 ;
        RECT 103.305 216.455 103.525 216.735 ;
        RECT 104.005 216.565 104.245 216.965 ;
        RECT 102.965 216.115 103.370 216.285 ;
        RECT 103.705 216.195 104.245 216.565 ;
        RECT 104.415 216.780 104.735 217.135 ;
        RECT 104.980 217.055 105.285 217.515 ;
        RECT 105.455 216.805 105.710 217.335 ;
        RECT 104.415 216.605 104.740 216.780 ;
        RECT 104.415 216.305 105.330 216.605 ;
        RECT 104.590 216.275 105.330 216.305 ;
        RECT 102.065 215.945 102.740 216.105 ;
        RECT 103.200 216.025 103.370 216.115 ;
        RECT 102.065 215.935 103.030 215.945 ;
        RECT 101.705 215.765 101.875 215.905 ;
        RECT 98.450 214.965 98.700 215.425 ;
        RECT 98.870 215.135 99.120 215.465 ;
        RECT 99.335 215.135 100.015 215.465 ;
        RECT 100.185 215.565 101.260 215.735 ;
        RECT 101.705 215.595 102.265 215.765 ;
        RECT 102.570 215.645 103.030 215.935 ;
        RECT 103.200 215.855 104.420 216.025 ;
        RECT 100.185 215.225 100.355 215.565 ;
        RECT 100.590 214.965 100.920 215.395 ;
        RECT 101.090 215.225 101.260 215.565 ;
        RECT 101.555 214.965 101.925 215.425 ;
        RECT 102.095 215.135 102.265 215.595 ;
        RECT 103.200 215.475 103.370 215.855 ;
        RECT 104.590 215.685 104.760 216.275 ;
        RECT 105.500 216.155 105.710 216.805 ;
        RECT 105.885 216.790 106.175 217.515 ;
        RECT 107.265 217.005 107.570 217.515 ;
        RECT 107.265 216.275 107.580 216.835 ;
        RECT 107.750 216.525 108.000 217.335 ;
        RECT 108.170 216.990 108.430 217.515 ;
        RECT 108.610 216.525 108.860 217.335 ;
        RECT 109.030 216.955 109.290 217.515 ;
        RECT 109.460 216.865 109.720 217.320 ;
        RECT 109.890 217.035 110.150 217.515 ;
        RECT 110.320 216.865 110.580 217.320 ;
        RECT 110.750 217.035 111.010 217.515 ;
        RECT 111.180 216.865 111.440 217.320 ;
        RECT 111.610 217.035 111.855 217.515 ;
        RECT 112.025 216.865 112.300 217.320 ;
        RECT 112.470 217.035 112.715 217.515 ;
        RECT 112.885 216.865 113.145 217.320 ;
        RECT 113.325 217.035 113.575 217.515 ;
        RECT 113.745 216.865 114.005 217.320 ;
        RECT 114.185 217.035 114.435 217.515 ;
        RECT 114.605 216.865 114.865 217.320 ;
        RECT 115.045 217.035 115.305 217.515 ;
        RECT 115.475 216.865 115.735 217.320 ;
        RECT 115.905 217.035 116.205 217.515 ;
        RECT 109.460 216.695 116.205 216.865 ;
        RECT 107.750 216.275 114.870 216.525 ;
        RECT 107.325 216.235 107.495 216.275 ;
        RECT 102.500 215.135 103.370 215.475 ;
        RECT 103.960 215.515 104.760 215.685 ;
        RECT 103.540 214.965 103.790 215.425 ;
        RECT 103.960 215.225 104.130 215.515 ;
        RECT 104.310 214.965 104.640 215.345 ;
        RECT 104.980 214.965 105.285 216.105 ;
        RECT 105.455 215.275 105.710 216.155 ;
        RECT 105.885 214.965 106.175 216.130 ;
        RECT 107.275 214.965 107.570 215.775 ;
        RECT 107.750 215.135 107.995 216.275 ;
        RECT 108.170 214.965 108.430 215.775 ;
        RECT 108.610 215.140 108.860 216.275 ;
        RECT 115.040 216.105 116.205 216.695 ;
        RECT 116.465 216.765 117.675 217.515 ;
        RECT 117.935 216.965 118.105 217.255 ;
        RECT 118.275 217.135 118.605 217.515 ;
        RECT 117.935 216.795 118.600 216.965 ;
        RECT 116.465 216.225 116.985 216.765 ;
        RECT 109.460 215.880 116.205 216.105 ;
        RECT 117.155 216.055 117.675 216.595 ;
        RECT 109.460 215.865 114.865 215.880 ;
        RECT 109.030 214.970 109.290 215.765 ;
        RECT 109.460 215.140 109.720 215.865 ;
        RECT 109.890 214.970 110.150 215.695 ;
        RECT 110.320 215.140 110.580 215.865 ;
        RECT 110.750 214.970 111.010 215.695 ;
        RECT 111.180 215.140 111.440 215.865 ;
        RECT 111.610 214.970 111.870 215.695 ;
        RECT 112.040 215.140 112.300 215.865 ;
        RECT 112.470 214.970 112.715 215.695 ;
        RECT 112.885 215.140 113.145 215.865 ;
        RECT 113.330 214.970 113.575 215.695 ;
        RECT 113.745 215.140 114.005 215.865 ;
        RECT 114.190 214.970 114.435 215.695 ;
        RECT 114.605 215.140 114.865 215.865 ;
        RECT 115.050 214.970 115.305 215.695 ;
        RECT 115.475 215.140 115.765 215.880 ;
        RECT 109.030 214.965 115.305 214.970 ;
        RECT 115.935 214.965 116.205 215.710 ;
        RECT 116.465 214.965 117.675 216.055 ;
        RECT 117.850 215.975 118.200 216.625 ;
        RECT 118.370 215.805 118.600 216.795 ;
        RECT 117.935 215.635 118.600 215.805 ;
        RECT 117.935 215.135 118.105 215.635 ;
        RECT 118.275 214.965 118.605 215.465 ;
        RECT 118.775 215.135 118.960 217.255 ;
        RECT 119.215 217.055 119.465 217.515 ;
        RECT 119.635 217.065 119.970 217.235 ;
        RECT 120.165 217.065 120.840 217.235 ;
        RECT 119.635 216.925 119.805 217.065 ;
        RECT 119.130 215.935 119.410 216.885 ;
        RECT 119.580 216.795 119.805 216.925 ;
        RECT 119.580 215.690 119.750 216.795 ;
        RECT 119.975 216.645 120.500 216.865 ;
        RECT 119.920 215.880 120.160 216.475 ;
        RECT 120.330 215.945 120.500 216.645 ;
        RECT 120.670 216.285 120.840 217.065 ;
        RECT 121.160 217.015 121.530 217.515 ;
        RECT 121.710 217.065 122.115 217.235 ;
        RECT 122.285 217.065 123.070 217.235 ;
        RECT 121.710 216.835 121.880 217.065 ;
        RECT 121.050 216.535 121.880 216.835 ;
        RECT 122.265 216.565 122.730 216.895 ;
        RECT 121.050 216.505 121.250 216.535 ;
        RECT 121.370 216.285 121.540 216.355 ;
        RECT 120.670 216.115 121.540 216.285 ;
        RECT 121.030 216.025 121.540 216.115 ;
        RECT 119.580 215.560 119.885 215.690 ;
        RECT 120.330 215.580 120.860 215.945 ;
        RECT 119.200 214.965 119.465 215.425 ;
        RECT 119.635 215.135 119.885 215.560 ;
        RECT 121.030 215.410 121.200 216.025 ;
        RECT 120.095 215.240 121.200 215.410 ;
        RECT 121.370 214.965 121.540 215.765 ;
        RECT 121.710 215.465 121.880 216.535 ;
        RECT 122.050 215.635 122.240 216.355 ;
        RECT 122.410 215.605 122.730 216.565 ;
        RECT 122.900 216.605 123.070 217.065 ;
        RECT 123.345 216.985 123.555 217.515 ;
        RECT 123.815 216.775 124.145 217.300 ;
        RECT 124.315 216.905 124.485 217.515 ;
        RECT 124.655 216.860 124.985 217.295 ;
        RECT 124.655 216.775 125.035 216.860 ;
        RECT 123.945 216.605 124.145 216.775 ;
        RECT 124.810 216.735 125.035 216.775 ;
        RECT 122.900 216.275 123.775 216.605 ;
        RECT 123.945 216.275 124.695 216.605 ;
        RECT 121.710 215.135 121.960 215.465 ;
        RECT 122.900 215.435 123.070 216.275 ;
        RECT 123.945 216.070 124.135 216.275 ;
        RECT 124.865 216.155 125.035 216.735 ;
        RECT 125.265 216.695 125.475 217.515 ;
        RECT 125.645 216.715 125.975 217.345 ;
        RECT 124.820 216.105 125.035 216.155 ;
        RECT 125.645 216.115 125.895 216.715 ;
        RECT 126.145 216.695 126.375 217.515 ;
        RECT 127.045 217.015 127.305 217.345 ;
        RECT 127.615 217.135 127.945 217.515 ;
        RECT 128.125 217.175 129.605 217.345 ;
        RECT 126.065 216.275 126.395 216.525 ;
        RECT 127.045 216.315 127.215 217.015 ;
        RECT 128.125 216.845 128.525 217.175 ;
        RECT 127.565 216.655 127.775 216.835 ;
        RECT 127.565 216.485 128.185 216.655 ;
        RECT 128.355 216.365 128.525 216.845 ;
        RECT 128.715 216.675 129.265 217.005 ;
        RECT 127.045 216.145 128.175 216.315 ;
        RECT 128.355 216.195 128.925 216.365 ;
        RECT 123.240 215.695 124.135 216.070 ;
        RECT 124.645 216.025 125.035 216.105 ;
        RECT 122.185 215.265 123.070 215.435 ;
        RECT 123.250 214.965 123.565 215.465 ;
        RECT 123.795 215.135 124.135 215.695 ;
        RECT 124.305 214.965 124.475 215.975 ;
        RECT 124.645 215.180 124.975 216.025 ;
        RECT 125.265 214.965 125.475 216.105 ;
        RECT 125.645 215.135 125.975 216.115 ;
        RECT 126.145 214.965 126.375 216.105 ;
        RECT 127.045 215.465 127.215 216.145 ;
        RECT 128.005 216.025 128.175 216.145 ;
        RECT 127.385 215.645 127.735 215.975 ;
        RECT 128.005 215.855 128.585 216.025 ;
        RECT 128.755 215.685 128.925 216.195 ;
        RECT 128.185 215.515 128.925 215.685 ;
        RECT 129.095 215.685 129.265 216.675 ;
        RECT 129.435 216.275 129.605 217.175 ;
        RECT 129.855 216.605 130.040 217.185 ;
        RECT 130.310 216.605 130.505 217.180 ;
        RECT 130.715 217.135 131.045 217.515 ;
        RECT 129.855 216.275 130.085 216.605 ;
        RECT 130.310 216.275 130.565 216.605 ;
        RECT 129.855 215.965 130.040 216.275 ;
        RECT 130.310 215.965 130.505 216.275 ;
        RECT 130.325 215.895 130.495 215.965 ;
        RECT 130.875 215.685 131.045 216.605 ;
        RECT 129.095 215.515 131.045 215.685 ;
        RECT 127.045 215.135 127.305 215.465 ;
        RECT 127.615 214.965 127.945 215.345 ;
        RECT 128.185 215.135 128.375 215.515 ;
        RECT 128.625 214.965 128.955 215.345 ;
        RECT 129.165 215.135 129.335 215.515 ;
        RECT 129.530 214.965 129.860 215.345 ;
        RECT 130.120 215.135 130.290 215.515 ;
        RECT 130.715 214.965 131.045 215.345 ;
        RECT 131.215 215.135 131.475 217.345 ;
        RECT 131.645 216.790 131.935 217.515 ;
        RECT 132.105 216.840 132.365 217.345 ;
        RECT 132.545 217.135 132.875 217.515 ;
        RECT 133.055 216.965 133.225 217.345 ;
        RECT 131.645 214.965 131.935 216.130 ;
        RECT 132.105 216.040 132.275 216.840 ;
        RECT 132.560 216.795 133.225 216.965 ;
        RECT 134.405 216.840 134.665 217.345 ;
        RECT 134.845 217.135 135.175 217.515 ;
        RECT 135.355 216.965 135.525 217.345 ;
        RECT 132.560 216.540 132.730 216.795 ;
        RECT 132.445 216.210 132.730 216.540 ;
        RECT 132.965 216.245 133.295 216.615 ;
        RECT 133.085 216.235 133.255 216.245 ;
        RECT 132.560 216.065 132.730 216.210 ;
        RECT 132.105 215.135 132.375 216.040 ;
        RECT 132.560 215.895 133.225 216.065 ;
        RECT 132.545 214.965 132.875 215.725 ;
        RECT 133.055 215.135 133.225 215.895 ;
        RECT 134.405 216.040 134.575 216.840 ;
        RECT 134.860 216.795 135.525 216.965 ;
        RECT 134.860 216.540 135.030 216.795 ;
        RECT 135.785 216.765 136.995 217.515 ;
        RECT 137.215 216.860 137.545 217.295 ;
        RECT 137.715 216.905 137.885 217.515 ;
        RECT 137.165 216.775 137.545 216.860 ;
        RECT 138.055 216.775 138.385 217.300 ;
        RECT 138.645 216.985 138.855 217.515 ;
        RECT 139.130 217.065 139.915 217.235 ;
        RECT 140.085 217.065 140.490 217.235 ;
        RECT 134.745 216.210 135.030 216.540 ;
        RECT 135.265 216.245 135.595 216.615 ;
        RECT 135.385 216.235 135.555 216.245 ;
        RECT 135.785 216.225 136.305 216.765 ;
        RECT 137.165 216.735 137.390 216.775 ;
        RECT 134.860 216.065 135.030 216.210 ;
        RECT 134.405 215.135 134.675 216.040 ;
        RECT 134.860 215.895 135.525 216.065 ;
        RECT 136.475 216.055 136.995 216.595 ;
        RECT 134.845 214.965 135.175 215.725 ;
        RECT 135.355 215.135 135.525 215.895 ;
        RECT 135.785 214.965 136.995 216.055 ;
        RECT 137.165 216.155 137.335 216.735 ;
        RECT 138.055 216.605 138.255 216.775 ;
        RECT 139.130 216.605 139.300 217.065 ;
        RECT 137.505 216.275 138.255 216.605 ;
        RECT 138.425 216.275 139.300 216.605 ;
        RECT 137.165 216.105 137.380 216.155 ;
        RECT 137.165 216.025 137.555 216.105 ;
        RECT 137.225 215.180 137.555 216.025 ;
        RECT 138.065 216.070 138.255 216.275 ;
        RECT 137.725 214.965 137.895 215.975 ;
        RECT 138.065 215.695 138.960 216.070 ;
        RECT 138.065 215.135 138.405 215.695 ;
        RECT 138.635 214.965 138.950 215.465 ;
        RECT 139.130 215.435 139.300 216.275 ;
        RECT 139.470 216.565 139.935 216.895 ;
        RECT 140.320 216.835 140.490 217.065 ;
        RECT 140.670 217.015 141.040 217.515 ;
        RECT 141.360 217.065 142.035 217.235 ;
        RECT 142.230 217.065 142.565 217.235 ;
        RECT 139.470 215.605 139.790 216.565 ;
        RECT 140.320 216.535 141.150 216.835 ;
        RECT 139.960 215.635 140.150 216.355 ;
        RECT 140.320 215.465 140.490 216.535 ;
        RECT 140.950 216.505 141.150 216.535 ;
        RECT 140.660 216.285 140.830 216.355 ;
        RECT 141.360 216.285 141.530 217.065 ;
        RECT 142.395 216.925 142.565 217.065 ;
        RECT 142.735 217.055 142.985 217.515 ;
        RECT 140.660 216.115 141.530 216.285 ;
        RECT 141.700 216.645 142.225 216.865 ;
        RECT 142.395 216.795 142.620 216.925 ;
        RECT 140.660 216.025 141.170 216.115 ;
        RECT 139.130 215.265 140.015 215.435 ;
        RECT 140.240 215.135 140.490 215.465 ;
        RECT 140.660 214.965 140.830 215.765 ;
        RECT 141.000 215.410 141.170 216.025 ;
        RECT 141.700 215.945 141.870 216.645 ;
        RECT 141.340 215.580 141.870 215.945 ;
        RECT 142.040 215.880 142.280 216.475 ;
        RECT 142.450 215.690 142.620 216.795 ;
        RECT 142.790 215.935 143.070 216.885 ;
        RECT 142.315 215.560 142.620 215.690 ;
        RECT 141.000 215.240 142.105 215.410 ;
        RECT 142.315 215.135 142.565 215.560 ;
        RECT 142.735 214.965 143.000 215.425 ;
        RECT 143.240 215.135 143.425 217.255 ;
        RECT 143.595 217.135 143.925 217.515 ;
        RECT 144.095 216.965 144.265 217.255 ;
        RECT 143.600 216.795 144.265 216.965 ;
        RECT 144.525 216.840 144.785 217.345 ;
        RECT 144.965 217.135 145.295 217.515 ;
        RECT 145.475 216.965 145.645 217.345 ;
        RECT 143.600 215.805 143.830 216.795 ;
        RECT 144.000 215.975 144.350 216.625 ;
        RECT 144.525 216.040 144.695 216.840 ;
        RECT 144.980 216.795 145.645 216.965 ;
        RECT 145.905 216.840 146.165 217.345 ;
        RECT 146.345 217.135 146.675 217.515 ;
        RECT 146.855 216.965 147.025 217.345 ;
        RECT 144.980 216.540 145.150 216.795 ;
        RECT 144.865 216.210 145.150 216.540 ;
        RECT 145.385 216.245 145.715 216.615 ;
        RECT 145.505 216.235 145.675 216.245 ;
        RECT 144.980 216.065 145.150 216.210 ;
        RECT 143.600 215.635 144.265 215.805 ;
        RECT 143.595 214.965 143.925 215.465 ;
        RECT 144.095 215.135 144.265 215.635 ;
        RECT 144.525 215.135 144.795 216.040 ;
        RECT 144.980 215.895 145.645 216.065 ;
        RECT 144.965 214.965 145.295 215.725 ;
        RECT 145.475 215.135 145.645 215.895 ;
        RECT 145.905 216.040 146.075 216.840 ;
        RECT 146.360 216.795 147.025 216.965 ;
        RECT 147.375 216.965 147.545 217.255 ;
        RECT 147.715 217.135 148.045 217.515 ;
        RECT 147.375 216.795 148.040 216.965 ;
        RECT 146.360 216.540 146.530 216.795 ;
        RECT 146.245 216.210 146.530 216.540 ;
        RECT 146.765 216.245 147.095 216.615 ;
        RECT 146.885 216.235 147.055 216.245 ;
        RECT 146.360 216.065 146.530 216.210 ;
        RECT 145.905 215.135 146.175 216.040 ;
        RECT 146.360 215.895 147.025 216.065 ;
        RECT 147.290 215.975 147.640 216.625 ;
        RECT 146.345 214.965 146.675 215.725 ;
        RECT 146.855 215.135 147.025 215.895 ;
        RECT 147.810 215.805 148.040 216.795 ;
        RECT 147.375 215.635 148.040 215.805 ;
        RECT 147.375 215.135 147.545 215.635 ;
        RECT 147.715 214.965 148.045 215.465 ;
        RECT 148.215 215.135 148.400 217.255 ;
        RECT 148.655 217.055 148.905 217.515 ;
        RECT 149.075 217.065 149.410 217.235 ;
        RECT 149.605 217.065 150.280 217.235 ;
        RECT 149.075 216.925 149.245 217.065 ;
        RECT 148.570 215.935 148.850 216.885 ;
        RECT 149.020 216.795 149.245 216.925 ;
        RECT 149.020 215.690 149.190 216.795 ;
        RECT 149.415 216.645 149.940 216.865 ;
        RECT 149.360 215.880 149.600 216.475 ;
        RECT 149.770 215.945 149.940 216.645 ;
        RECT 150.110 216.285 150.280 217.065 ;
        RECT 150.600 217.015 150.970 217.515 ;
        RECT 151.150 217.065 151.555 217.235 ;
        RECT 151.725 217.065 152.510 217.235 ;
        RECT 151.150 216.835 151.320 217.065 ;
        RECT 150.490 216.535 151.320 216.835 ;
        RECT 151.705 216.565 152.170 216.895 ;
        RECT 150.490 216.505 150.690 216.535 ;
        RECT 150.810 216.285 150.980 216.355 ;
        RECT 150.110 216.115 150.980 216.285 ;
        RECT 150.470 216.025 150.980 216.115 ;
        RECT 149.020 215.560 149.325 215.690 ;
        RECT 149.770 215.580 150.300 215.945 ;
        RECT 148.640 214.965 148.905 215.425 ;
        RECT 149.075 215.135 149.325 215.560 ;
        RECT 150.470 215.410 150.640 216.025 ;
        RECT 149.535 215.240 150.640 215.410 ;
        RECT 150.810 214.965 150.980 215.765 ;
        RECT 151.150 215.465 151.320 216.535 ;
        RECT 151.490 215.635 151.680 216.355 ;
        RECT 151.850 215.605 152.170 216.565 ;
        RECT 152.340 216.605 152.510 217.065 ;
        RECT 152.785 216.985 152.995 217.515 ;
        RECT 153.255 216.775 153.585 217.300 ;
        RECT 153.755 216.905 153.925 217.515 ;
        RECT 154.095 216.860 154.425 217.295 ;
        RECT 154.095 216.775 154.475 216.860 ;
        RECT 153.385 216.605 153.585 216.775 ;
        RECT 154.250 216.735 154.475 216.775 ;
        RECT 152.340 216.275 153.215 216.605 ;
        RECT 153.385 216.275 154.135 216.605 ;
        RECT 151.150 215.135 151.400 215.465 ;
        RECT 152.340 215.435 152.510 216.275 ;
        RECT 153.385 216.070 153.575 216.275 ;
        RECT 154.305 216.155 154.475 216.735 ;
        RECT 154.260 216.105 154.475 216.155 ;
        RECT 152.680 215.695 153.575 216.070 ;
        RECT 154.085 216.025 154.475 216.105 ;
        RECT 154.645 216.840 154.905 217.345 ;
        RECT 155.085 217.135 155.415 217.515 ;
        RECT 155.595 216.965 155.765 217.345 ;
        RECT 154.645 216.040 154.815 216.840 ;
        RECT 155.100 216.795 155.765 216.965 ;
        RECT 155.100 216.540 155.270 216.795 ;
        RECT 156.945 216.765 158.155 217.515 ;
        RECT 154.985 216.210 155.270 216.540 ;
        RECT 155.505 216.245 155.835 216.615 ;
        RECT 155.625 216.235 155.795 216.245 ;
        RECT 155.100 216.065 155.270 216.210 ;
        RECT 151.625 215.265 152.510 215.435 ;
        RECT 152.690 214.965 153.005 215.465 ;
        RECT 153.235 215.135 153.575 215.695 ;
        RECT 153.745 214.965 153.915 215.975 ;
        RECT 154.085 215.180 154.415 216.025 ;
        RECT 154.645 215.135 154.915 216.040 ;
        RECT 155.100 215.895 155.765 216.065 ;
        RECT 155.085 214.965 155.415 215.725 ;
        RECT 155.595 215.135 155.765 215.895 ;
        RECT 156.945 216.055 157.465 216.595 ;
        RECT 157.635 216.225 158.155 216.765 ;
        RECT 156.945 214.965 158.155 216.055 ;
        RECT 2.760 214.795 158.240 214.965 ;
        RECT 2.845 213.705 4.055 214.795 ;
        RECT 4.225 214.360 9.570 214.795 ;
        RECT 9.745 214.360 15.090 214.795 ;
        RECT 2.845 212.995 3.365 213.535 ;
        RECT 3.535 213.165 4.055 213.705 ;
        RECT 2.845 212.245 4.055 212.995 ;
        RECT 5.810 212.790 6.150 213.620 ;
        RECT 7.630 213.110 7.980 214.360 ;
        RECT 11.330 212.790 11.670 213.620 ;
        RECT 13.150 213.110 13.500 214.360 ;
        RECT 15.725 213.630 16.015 214.795 ;
        RECT 16.185 214.360 21.530 214.795 ;
        RECT 21.705 214.360 27.050 214.795 ;
        RECT 27.225 214.360 32.570 214.795 ;
        RECT 32.745 214.360 38.090 214.795 ;
        RECT 4.225 212.245 9.570 212.790 ;
        RECT 9.745 212.245 15.090 212.790 ;
        RECT 15.725 212.245 16.015 212.970 ;
        RECT 17.770 212.790 18.110 213.620 ;
        RECT 19.590 213.110 19.940 214.360 ;
        RECT 23.290 212.790 23.630 213.620 ;
        RECT 25.110 213.110 25.460 214.360 ;
        RECT 28.810 212.790 29.150 213.620 ;
        RECT 30.630 213.110 30.980 214.360 ;
        RECT 34.330 212.790 34.670 213.620 ;
        RECT 36.150 213.110 36.500 214.360 ;
        RECT 38.265 213.705 40.855 214.795 ;
        RECT 38.265 213.015 39.475 213.535 ;
        RECT 39.645 213.185 40.855 213.705 ;
        RECT 41.485 213.630 41.775 214.795 ;
        RECT 41.945 214.360 47.290 214.795 ;
        RECT 47.465 214.360 52.810 214.795 ;
        RECT 16.185 212.245 21.530 212.790 ;
        RECT 21.705 212.245 27.050 212.790 ;
        RECT 27.225 212.245 32.570 212.790 ;
        RECT 32.745 212.245 38.090 212.790 ;
        RECT 38.265 212.245 40.855 213.015 ;
        RECT 41.485 212.245 41.775 212.970 ;
        RECT 43.530 212.790 43.870 213.620 ;
        RECT 45.350 213.110 45.700 214.360 ;
        RECT 49.050 212.790 49.390 213.620 ;
        RECT 50.870 213.110 51.220 214.360 ;
        RECT 52.985 213.705 54.195 214.795 ;
        RECT 54.420 213.925 54.705 214.795 ;
        RECT 54.875 214.165 55.135 214.625 ;
        RECT 55.310 214.335 55.565 214.795 ;
        RECT 55.735 214.165 55.995 214.625 ;
        RECT 54.875 213.995 55.995 214.165 ;
        RECT 56.165 213.995 56.475 214.795 ;
        RECT 54.875 213.745 55.135 213.995 ;
        RECT 56.645 213.825 56.955 214.625 ;
        RECT 57.180 213.925 57.465 214.795 ;
        RECT 57.635 214.165 57.895 214.625 ;
        RECT 58.070 214.335 58.325 214.795 ;
        RECT 58.495 214.165 58.755 214.625 ;
        RECT 57.635 213.995 58.755 214.165 ;
        RECT 58.925 213.995 59.235 214.795 ;
        RECT 52.985 212.995 53.505 213.535 ;
        RECT 53.675 213.165 54.195 213.705 ;
        RECT 54.380 213.575 55.135 213.745 ;
        RECT 55.925 213.655 56.955 213.825 ;
        RECT 57.635 213.745 57.895 213.995 ;
        RECT 59.405 213.825 59.715 214.625 ;
        RECT 54.380 213.065 54.785 213.575 ;
        RECT 55.925 213.405 56.095 213.655 ;
        RECT 54.955 213.235 56.095 213.405 ;
        RECT 41.945 212.245 47.290 212.790 ;
        RECT 47.465 212.245 52.810 212.790 ;
        RECT 52.985 212.245 54.195 212.995 ;
        RECT 54.380 212.895 56.030 213.065 ;
        RECT 56.265 212.915 56.615 213.485 ;
        RECT 54.425 212.245 54.705 212.725 ;
        RECT 54.875 212.505 55.135 212.895 ;
        RECT 55.310 212.245 55.565 212.725 ;
        RECT 55.735 212.505 56.030 212.895 ;
        RECT 56.785 212.745 56.955 213.655 ;
        RECT 57.140 213.575 57.895 213.745 ;
        RECT 58.685 213.655 59.715 213.825 ;
        RECT 57.140 213.065 57.545 213.575 ;
        RECT 58.685 213.405 58.855 213.655 ;
        RECT 57.715 213.235 58.855 213.405 ;
        RECT 57.140 212.895 58.790 213.065 ;
        RECT 59.025 212.915 59.375 213.485 ;
        RECT 56.210 212.245 56.485 212.725 ;
        RECT 56.655 212.415 56.955 212.745 ;
        RECT 57.185 212.245 57.465 212.725 ;
        RECT 57.635 212.505 57.895 212.895 ;
        RECT 58.070 212.245 58.325 212.725 ;
        RECT 58.495 212.505 58.790 212.895 ;
        RECT 59.545 212.745 59.715 213.655 ;
        RECT 58.970 212.245 59.245 212.725 ;
        RECT 59.415 212.415 59.715 212.745 ;
        RECT 59.885 212.415 60.145 214.625 ;
        RECT 60.315 214.415 60.645 214.795 ;
        RECT 61.070 214.245 61.240 214.625 ;
        RECT 61.500 214.415 61.830 214.795 ;
        RECT 62.025 214.245 62.195 214.625 ;
        RECT 62.405 214.415 62.735 214.795 ;
        RECT 62.985 214.245 63.175 214.625 ;
        RECT 63.415 214.415 63.745 214.795 ;
        RECT 64.055 214.295 64.315 214.625 ;
        RECT 60.315 214.075 62.265 214.245 ;
        RECT 60.315 213.155 60.485 214.075 ;
        RECT 60.855 213.485 61.050 213.795 ;
        RECT 61.320 213.485 61.505 213.795 ;
        RECT 60.795 213.155 61.050 213.485 ;
        RECT 61.275 213.155 61.505 213.485 ;
        RECT 60.315 212.245 60.645 212.625 ;
        RECT 60.855 212.580 61.050 213.155 ;
        RECT 61.320 212.575 61.505 213.155 ;
        RECT 61.755 212.585 61.925 213.485 ;
        RECT 62.095 213.085 62.265 214.075 ;
        RECT 62.435 214.075 63.175 214.245 ;
        RECT 62.435 213.565 62.605 214.075 ;
        RECT 62.775 213.735 63.355 213.905 ;
        RECT 63.625 213.785 63.975 214.115 ;
        RECT 63.185 213.615 63.355 213.735 ;
        RECT 64.145 213.615 64.315 214.295 ;
        RECT 62.435 213.395 63.005 213.565 ;
        RECT 63.185 213.445 64.315 213.615 ;
        RECT 62.095 212.755 62.645 213.085 ;
        RECT 62.835 212.915 63.005 213.395 ;
        RECT 63.175 213.105 63.795 213.275 ;
        RECT 63.585 212.925 63.795 213.105 ;
        RECT 62.835 212.585 63.235 212.915 ;
        RECT 64.145 212.745 64.315 213.445 ;
        RECT 61.755 212.415 63.235 212.585 ;
        RECT 63.415 212.245 63.745 212.625 ;
        RECT 64.055 212.415 64.315 212.745 ;
        RECT 64.485 213.825 64.795 214.625 ;
        RECT 64.965 213.995 65.275 214.795 ;
        RECT 65.445 214.165 65.705 214.625 ;
        RECT 65.875 214.335 66.130 214.795 ;
        RECT 66.305 214.165 66.565 214.625 ;
        RECT 65.445 213.995 66.565 214.165 ;
        RECT 64.485 213.655 65.515 213.825 ;
        RECT 64.485 212.745 64.655 213.655 ;
        RECT 64.825 212.915 65.175 213.485 ;
        RECT 65.345 213.405 65.515 213.655 ;
        RECT 66.305 213.745 66.565 213.995 ;
        RECT 66.735 213.925 67.020 214.795 ;
        RECT 66.305 213.575 67.060 213.745 ;
        RECT 67.245 213.630 67.535 214.795 ;
        RECT 67.870 214.455 69.965 214.625 ;
        RECT 67.870 214.075 68.285 214.455 ;
        RECT 68.455 213.905 68.625 214.285 ;
        RECT 68.795 214.095 69.125 214.455 ;
        RECT 69.295 213.905 69.465 214.285 ;
        RECT 65.345 213.235 66.485 213.405 ;
        RECT 66.655 213.065 67.060 213.575 ;
        RECT 65.410 212.895 67.060 213.065 ;
        RECT 67.705 213.605 69.465 213.905 ;
        RECT 69.635 213.825 69.965 214.455 ;
        RECT 70.135 213.995 70.385 214.795 ;
        RECT 70.555 213.825 70.725 214.625 ;
        RECT 70.895 213.995 71.225 214.795 ;
        RECT 71.395 213.825 71.670 214.625 ;
        RECT 69.635 213.615 71.670 213.825 ;
        RECT 71.845 213.705 73.515 214.795 ;
        RECT 73.685 214.200 73.945 214.380 ;
        RECT 74.150 214.370 74.510 214.795 ;
        RECT 75.020 214.370 75.350 214.795 ;
        RECT 75.855 214.370 76.195 214.795 ;
        RECT 77.120 214.370 77.655 214.585 ;
        RECT 73.685 214.030 77.220 214.200 ;
        RECT 73.685 213.970 74.365 214.030 ;
        RECT 67.705 213.065 68.105 213.605 ;
        RECT 68.275 213.235 69.640 213.435 ;
        RECT 69.960 213.235 71.620 213.435 ;
        RECT 64.485 212.415 64.785 212.745 ;
        RECT 64.955 212.245 65.230 212.725 ;
        RECT 65.410 212.505 65.705 212.895 ;
        RECT 65.875 212.245 66.130 212.725 ;
        RECT 66.305 212.505 66.565 212.895 ;
        RECT 66.735 212.245 67.015 212.725 ;
        RECT 67.245 212.245 67.535 212.970 ;
        RECT 67.705 212.885 71.225 213.065 ;
        RECT 67.920 212.245 68.205 212.715 ;
        RECT 68.375 212.415 68.705 212.885 ;
        RECT 68.875 212.245 69.045 212.715 ;
        RECT 69.215 212.415 69.545 212.885 ;
        RECT 69.715 212.245 69.885 212.715 ;
        RECT 70.055 212.415 70.385 212.885 ;
        RECT 70.555 212.245 70.725 212.715 ;
        RECT 70.895 212.415 71.225 212.885 ;
        RECT 71.395 212.245 71.670 213.065 ;
        RECT 71.845 213.015 72.595 213.535 ;
        RECT 72.765 213.185 73.515 213.705 ;
        RECT 73.685 213.235 74.025 213.800 ;
        RECT 74.195 213.065 74.365 213.970 ;
        RECT 71.845 212.245 73.515 213.015 ;
        RECT 73.685 212.895 74.365 213.065 ;
        RECT 74.535 213.575 75.820 213.860 ;
        RECT 76.000 213.575 76.320 213.860 ;
        RECT 74.535 213.065 74.705 213.575 ;
        RECT 74.875 213.235 75.965 213.405 ;
        RECT 74.535 212.895 75.625 213.065 ;
        RECT 73.685 212.450 73.945 212.895 ;
        RECT 74.220 212.245 74.390 212.725 ;
        RECT 74.600 212.445 74.930 212.895 ;
        RECT 75.455 212.745 75.625 212.895 ;
        RECT 75.795 213.050 75.965 213.235 ;
        RECT 76.135 213.155 76.320 213.575 ;
        RECT 76.490 213.155 76.800 213.860 ;
        RECT 76.990 213.485 77.220 214.030 ;
        RECT 76.990 213.155 77.280 213.485 ;
        RECT 75.795 212.985 76.000 213.050 ;
        RECT 77.450 212.985 77.655 214.370 ;
        RECT 77.990 214.455 80.085 214.625 ;
        RECT 77.990 214.075 78.405 214.455 ;
        RECT 78.575 213.905 78.745 214.285 ;
        RECT 78.915 214.095 79.245 214.455 ;
        RECT 79.415 213.905 79.585 214.285 ;
        RECT 75.795 212.880 77.655 212.985 ;
        RECT 77.825 213.605 79.585 213.905 ;
        RECT 79.755 213.825 80.085 214.455 ;
        RECT 80.255 213.995 80.505 214.795 ;
        RECT 80.675 213.825 80.845 214.625 ;
        RECT 81.015 213.995 81.345 214.795 ;
        RECT 81.515 213.825 81.790 214.625 ;
        RECT 82.055 214.050 82.325 214.795 ;
        RECT 82.955 214.790 89.230 214.795 ;
        RECT 82.495 213.880 82.785 214.620 ;
        RECT 82.955 214.065 83.210 214.790 ;
        RECT 83.395 213.895 83.655 214.620 ;
        RECT 83.825 214.065 84.070 214.790 ;
        RECT 84.255 213.895 84.515 214.620 ;
        RECT 84.685 214.065 84.930 214.790 ;
        RECT 85.115 213.895 85.375 214.620 ;
        RECT 85.545 214.065 85.790 214.790 ;
        RECT 85.960 213.895 86.220 214.620 ;
        RECT 86.390 214.065 86.650 214.790 ;
        RECT 86.820 213.895 87.080 214.620 ;
        RECT 87.250 214.065 87.510 214.790 ;
        RECT 87.680 213.895 87.940 214.620 ;
        RECT 88.110 214.065 88.370 214.790 ;
        RECT 88.540 213.895 88.800 214.620 ;
        RECT 88.970 213.995 89.230 214.790 ;
        RECT 83.395 213.880 88.800 213.895 ;
        RECT 79.755 213.615 81.790 213.825 ;
        RECT 82.055 213.655 88.800 213.880 ;
        RECT 77.825 213.065 78.225 213.605 ;
        RECT 78.395 213.235 79.760 213.435 ;
        RECT 80.080 213.235 81.740 213.435 ;
        RECT 82.055 213.065 83.220 213.655 ;
        RECT 89.400 213.485 89.650 214.620 ;
        RECT 89.830 213.985 90.090 214.795 ;
        RECT 90.265 213.485 90.510 214.625 ;
        RECT 90.690 213.985 90.985 214.795 ;
        RECT 91.170 214.370 91.505 214.795 ;
        RECT 91.675 214.190 91.860 214.595 ;
        RECT 91.195 214.015 91.860 214.190 ;
        RECT 92.065 214.015 92.395 214.795 ;
        RECT 83.390 213.235 90.510 213.485 ;
        RECT 77.825 212.885 81.345 213.065 ;
        RECT 75.850 212.815 77.655 212.880 ;
        RECT 75.100 212.245 75.270 212.725 ;
        RECT 75.455 212.415 75.690 212.745 ;
        RECT 75.860 212.245 76.190 212.645 ;
        RECT 76.360 212.465 76.530 212.815 ;
        RECT 77.260 212.765 77.655 212.815 ;
        RECT 76.700 212.245 77.090 212.645 ;
        RECT 77.260 212.465 77.515 212.765 ;
        RECT 78.040 212.245 78.325 212.715 ;
        RECT 78.495 212.415 78.825 212.885 ;
        RECT 78.995 212.245 79.165 212.715 ;
        RECT 79.335 212.415 79.665 212.885 ;
        RECT 79.835 212.245 80.005 212.715 ;
        RECT 80.175 212.415 80.505 212.885 ;
        RECT 80.675 212.245 80.845 212.715 ;
        RECT 81.015 212.415 81.345 212.885 ;
        RECT 81.515 212.245 81.790 213.065 ;
        RECT 82.055 212.895 88.800 213.065 ;
        RECT 82.055 212.245 82.355 212.725 ;
        RECT 82.525 212.440 82.785 212.895 ;
        RECT 82.955 212.245 83.215 212.725 ;
        RECT 83.395 212.440 83.655 212.895 ;
        RECT 83.825 212.245 84.075 212.725 ;
        RECT 84.255 212.440 84.515 212.895 ;
        RECT 84.685 212.245 84.935 212.725 ;
        RECT 85.115 212.440 85.375 212.895 ;
        RECT 85.545 212.245 85.790 212.725 ;
        RECT 85.960 212.440 86.235 212.895 ;
        RECT 86.405 212.245 86.650 212.725 ;
        RECT 86.820 212.440 87.080 212.895 ;
        RECT 87.250 212.245 87.510 212.725 ;
        RECT 87.680 212.440 87.940 212.895 ;
        RECT 88.110 212.245 88.370 212.725 ;
        RECT 88.540 212.440 88.800 212.895 ;
        RECT 88.970 212.245 89.230 212.805 ;
        RECT 89.400 212.425 89.650 213.235 ;
        RECT 89.830 212.245 90.090 212.770 ;
        RECT 90.260 212.425 90.510 213.235 ;
        RECT 90.680 212.925 90.995 213.485 ;
        RECT 91.195 212.985 91.535 214.015 ;
        RECT 92.565 213.825 92.835 214.595 ;
        RECT 91.705 213.655 92.835 213.825 ;
        RECT 91.705 213.155 91.955 213.655 ;
        RECT 91.195 212.815 91.880 212.985 ;
        RECT 92.135 212.905 92.495 213.485 ;
        RECT 90.690 212.245 90.995 212.755 ;
        RECT 91.170 212.245 91.505 212.645 ;
        RECT 91.675 212.415 91.880 212.815 ;
        RECT 92.665 212.745 92.835 213.655 ;
        RECT 93.005 213.630 93.295 214.795 ;
        RECT 93.465 214.360 98.810 214.795 ;
        RECT 92.090 212.245 92.365 212.725 ;
        RECT 92.575 212.415 92.835 212.745 ;
        RECT 93.005 212.245 93.295 212.970 ;
        RECT 95.050 212.790 95.390 213.620 ;
        RECT 96.870 213.110 97.220 214.360 ;
        RECT 98.985 213.705 101.575 214.795 ;
        RECT 98.985 213.015 100.195 213.535 ;
        RECT 100.365 213.185 101.575 213.705 ;
        RECT 102.210 213.655 102.545 214.625 ;
        RECT 102.715 213.655 102.885 214.795 ;
        RECT 103.055 214.455 105.085 214.625 ;
        RECT 93.465 212.245 98.810 212.790 ;
        RECT 98.985 212.245 101.575 213.015 ;
        RECT 102.210 213.005 102.380 213.655 ;
        RECT 103.055 213.485 103.225 214.455 ;
        RECT 102.550 213.155 102.805 213.485 ;
        RECT 103.030 213.155 103.225 213.485 ;
        RECT 103.395 214.115 104.520 214.285 ;
        RECT 102.210 212.985 102.435 213.005 ;
        RECT 102.635 212.985 102.805 213.155 ;
        RECT 103.395 212.985 103.565 214.115 ;
        RECT 102.210 212.415 102.465 212.985 ;
        RECT 102.635 212.815 103.565 212.985 ;
        RECT 103.735 213.775 104.745 213.945 ;
        RECT 103.735 212.975 103.905 213.775 ;
        RECT 104.110 213.005 104.385 213.575 ;
        RECT 104.105 212.835 104.385 213.005 ;
        RECT 103.390 212.780 103.565 212.815 ;
        RECT 102.635 212.245 102.965 212.645 ;
        RECT 103.390 212.415 103.920 212.780 ;
        RECT 104.110 212.415 104.385 212.835 ;
        RECT 104.555 212.415 104.745 213.775 ;
        RECT 104.915 213.790 105.085 214.455 ;
        RECT 105.255 214.035 105.425 214.795 ;
        RECT 105.660 214.035 106.175 214.445 ;
        RECT 104.915 213.600 105.665 213.790 ;
        RECT 105.025 213.515 105.195 213.600 ;
        RECT 105.835 213.225 106.175 214.035 ;
        RECT 104.945 213.055 106.175 213.225 ;
        RECT 106.345 213.655 106.730 214.625 ;
        RECT 106.900 214.335 107.225 214.795 ;
        RECT 107.745 214.165 108.025 214.625 ;
        RECT 106.900 213.945 108.025 214.165 ;
        RECT 104.925 212.245 105.435 212.780 ;
        RECT 105.655 212.450 105.900 213.055 ;
        RECT 106.345 212.985 106.625 213.655 ;
        RECT 106.900 213.485 107.350 213.945 ;
        RECT 108.215 213.775 108.615 214.625 ;
        RECT 109.015 214.335 109.285 214.795 ;
        RECT 109.455 214.165 109.740 214.625 ;
        RECT 106.795 213.155 107.350 213.485 ;
        RECT 107.520 213.215 108.615 213.775 ;
        RECT 106.900 213.045 107.350 213.155 ;
        RECT 106.345 212.415 106.730 212.985 ;
        RECT 106.900 212.875 108.025 213.045 ;
        RECT 106.900 212.245 107.225 212.705 ;
        RECT 107.745 212.415 108.025 212.875 ;
        RECT 108.215 212.415 108.615 213.215 ;
        RECT 108.785 213.945 109.740 214.165 ;
        RECT 108.785 213.045 108.995 213.945 ;
        RECT 109.165 213.215 109.855 213.775 ;
        RECT 110.025 213.655 110.410 214.625 ;
        RECT 110.580 214.335 110.905 214.795 ;
        RECT 111.425 214.165 111.705 214.625 ;
        RECT 110.580 213.945 111.705 214.165 ;
        RECT 108.785 212.875 109.740 213.045 ;
        RECT 109.015 212.245 109.285 212.705 ;
        RECT 109.455 212.415 109.740 212.875 ;
        RECT 110.025 212.985 110.305 213.655 ;
        RECT 110.580 213.485 111.030 213.945 ;
        RECT 111.895 213.775 112.295 214.625 ;
        RECT 112.695 214.335 112.965 214.795 ;
        RECT 113.135 214.165 113.420 214.625 ;
        RECT 110.475 213.155 111.030 213.485 ;
        RECT 111.200 213.215 112.295 213.775 ;
        RECT 110.580 213.045 111.030 213.155 ;
        RECT 110.025 212.415 110.410 212.985 ;
        RECT 110.580 212.875 111.705 213.045 ;
        RECT 110.580 212.245 110.905 212.705 ;
        RECT 111.425 212.415 111.705 212.875 ;
        RECT 111.895 212.415 112.295 213.215 ;
        RECT 112.465 213.945 113.420 214.165 ;
        RECT 113.725 214.205 113.965 214.595 ;
        RECT 114.135 214.385 114.485 214.795 ;
        RECT 113.725 214.005 114.475 214.205 ;
        RECT 112.465 213.045 112.675 213.945 ;
        RECT 112.845 213.215 113.535 213.775 ;
        RECT 112.465 212.875 113.420 213.045 ;
        RECT 112.695 212.245 112.965 212.705 ;
        RECT 113.135 212.415 113.420 212.875 ;
        RECT 113.725 212.485 113.955 213.825 ;
        RECT 114.135 213.325 114.475 214.005 ;
        RECT 114.655 213.505 114.985 214.615 ;
        RECT 115.155 214.145 115.335 214.615 ;
        RECT 115.505 214.315 115.835 214.795 ;
        RECT 116.010 214.145 116.180 214.615 ;
        RECT 115.155 213.945 116.180 214.145 ;
        RECT 114.135 212.425 114.365 213.325 ;
        RECT 114.655 213.205 115.200 213.505 ;
        RECT 114.565 212.245 114.810 213.025 ;
        RECT 114.980 212.975 115.200 213.205 ;
        RECT 115.370 213.155 115.795 213.775 ;
        RECT 115.990 213.155 116.250 213.775 ;
        RECT 116.445 213.655 116.730 214.795 ;
        RECT 116.460 212.975 116.720 213.485 ;
        RECT 114.980 212.785 116.720 212.975 ;
        RECT 114.980 212.425 115.410 212.785 ;
        RECT 115.990 212.245 116.720 212.615 ;
        RECT 116.920 212.425 117.200 214.615 ;
        RECT 117.385 213.720 117.655 214.625 ;
        RECT 117.825 214.035 118.155 214.795 ;
        RECT 118.335 213.865 118.505 214.625 ;
        RECT 117.385 213.005 117.555 213.720 ;
        RECT 117.840 213.695 118.505 213.865 ;
        RECT 117.840 213.550 118.010 213.695 ;
        RECT 118.765 213.630 119.055 214.795 ;
        RECT 119.245 213.740 119.550 214.525 ;
        RECT 119.730 214.325 120.415 214.795 ;
        RECT 119.725 213.805 120.420 214.115 ;
        RECT 117.725 213.220 118.010 213.550 ;
        RECT 117.385 212.920 117.615 213.005 ;
        RECT 117.840 212.965 118.010 213.220 ;
        RECT 118.245 213.145 118.575 213.515 ;
        RECT 119.245 213.005 119.420 213.740 ;
        RECT 120.595 213.635 120.880 214.580 ;
        RECT 121.055 214.345 121.385 214.795 ;
        RECT 121.555 214.175 121.725 214.605 ;
        RECT 120.020 213.485 120.880 213.635 ;
        RECT 119.595 213.465 120.880 213.485 ;
        RECT 121.050 213.945 121.725 214.175 ;
        RECT 122.075 214.125 122.245 214.625 ;
        RECT 122.415 214.295 122.745 214.795 ;
        RECT 122.075 213.955 122.740 214.125 ;
        RECT 119.595 213.105 120.580 213.465 ;
        RECT 121.050 213.295 121.285 213.945 ;
        RECT 117.385 212.415 117.645 212.920 ;
        RECT 117.840 212.795 118.505 212.965 ;
        RECT 117.825 212.245 118.155 212.625 ;
        RECT 118.335 212.415 118.505 212.795 ;
        RECT 118.765 212.245 119.055 212.970 ;
        RECT 119.245 212.935 119.455 213.005 ;
        RECT 119.245 212.415 119.485 212.935 ;
        RECT 120.410 212.770 120.580 213.105 ;
        RECT 120.750 212.965 121.285 213.295 ;
        RECT 121.065 212.815 121.285 212.965 ;
        RECT 121.455 212.925 121.755 213.775 ;
        RECT 121.990 213.135 122.340 213.785 ;
        RECT 122.510 212.965 122.740 213.955 ;
        RECT 119.655 212.245 120.050 212.740 ;
        RECT 120.410 212.575 120.785 212.770 ;
        RECT 120.615 212.430 120.785 212.575 ;
        RECT 121.065 212.440 121.305 212.815 ;
        RECT 122.075 212.795 122.740 212.965 ;
        RECT 121.475 212.245 121.810 212.750 ;
        RECT 122.075 212.505 122.245 212.795 ;
        RECT 122.415 212.245 122.745 212.625 ;
        RECT 122.915 212.505 123.100 214.625 ;
        RECT 123.340 214.335 123.605 214.795 ;
        RECT 123.775 214.200 124.025 214.625 ;
        RECT 124.235 214.350 125.340 214.520 ;
        RECT 123.720 214.070 124.025 214.200 ;
        RECT 123.270 212.875 123.550 213.825 ;
        RECT 123.720 212.965 123.890 214.070 ;
        RECT 124.060 213.285 124.300 213.880 ;
        RECT 124.470 213.815 125.000 214.180 ;
        RECT 124.470 213.115 124.640 213.815 ;
        RECT 125.170 213.735 125.340 214.350 ;
        RECT 125.510 213.995 125.680 214.795 ;
        RECT 125.850 214.295 126.100 214.625 ;
        RECT 126.325 214.325 127.210 214.495 ;
        RECT 125.170 213.645 125.680 213.735 ;
        RECT 123.720 212.835 123.945 212.965 ;
        RECT 124.115 212.895 124.640 213.115 ;
        RECT 124.810 213.475 125.680 213.645 ;
        RECT 123.355 212.245 123.605 212.705 ;
        RECT 123.775 212.695 123.945 212.835 ;
        RECT 124.810 212.695 124.980 213.475 ;
        RECT 125.510 213.405 125.680 213.475 ;
        RECT 125.190 213.225 125.390 213.255 ;
        RECT 125.850 213.225 126.020 214.295 ;
        RECT 126.190 213.405 126.380 214.125 ;
        RECT 125.190 212.925 126.020 213.225 ;
        RECT 126.550 213.195 126.870 214.155 ;
        RECT 123.775 212.525 124.110 212.695 ;
        RECT 124.305 212.525 124.980 212.695 ;
        RECT 125.300 212.245 125.670 212.745 ;
        RECT 125.850 212.695 126.020 212.925 ;
        RECT 126.405 212.865 126.870 213.195 ;
        RECT 127.040 213.485 127.210 214.325 ;
        RECT 127.390 214.295 127.705 214.795 ;
        RECT 127.935 214.065 128.275 214.625 ;
        RECT 127.380 213.690 128.275 214.065 ;
        RECT 128.445 213.785 128.615 214.795 ;
        RECT 128.085 213.485 128.275 213.690 ;
        RECT 128.785 213.735 129.115 214.580 ;
        RECT 128.785 213.655 129.175 213.735 ;
        RECT 128.960 213.605 129.175 213.655 ;
        RECT 127.040 213.155 127.915 213.485 ;
        RECT 128.085 213.155 128.835 213.485 ;
        RECT 127.040 212.695 127.210 213.155 ;
        RECT 128.085 212.985 128.285 213.155 ;
        RECT 129.005 213.025 129.175 213.605 ;
        RECT 128.950 213.005 129.175 213.025 ;
        RECT 128.945 212.985 129.175 213.005 ;
        RECT 125.850 212.525 126.255 212.695 ;
        RECT 126.425 212.525 127.210 212.695 ;
        RECT 127.485 212.245 127.695 212.775 ;
        RECT 127.955 212.460 128.285 212.985 ;
        RECT 128.795 212.900 129.175 212.985 ;
        RECT 129.345 213.655 129.730 214.625 ;
        RECT 129.900 214.335 130.225 214.795 ;
        RECT 130.745 214.165 131.025 214.625 ;
        RECT 129.900 213.945 131.025 214.165 ;
        RECT 129.345 212.985 129.625 213.655 ;
        RECT 129.900 213.485 130.350 213.945 ;
        RECT 131.215 213.775 131.615 214.625 ;
        RECT 132.015 214.335 132.285 214.795 ;
        RECT 132.455 214.165 132.740 214.625 ;
        RECT 133.030 214.370 133.365 214.795 ;
        RECT 133.535 214.190 133.720 214.595 ;
        RECT 129.795 213.155 130.350 213.485 ;
        RECT 130.520 213.215 131.615 213.775 ;
        RECT 129.900 213.045 130.350 213.155 ;
        RECT 128.455 212.245 128.625 212.855 ;
        RECT 128.795 212.465 129.125 212.900 ;
        RECT 129.345 212.415 129.730 212.985 ;
        RECT 129.900 212.875 131.025 213.045 ;
        RECT 129.900 212.245 130.225 212.705 ;
        RECT 130.745 212.415 131.025 212.875 ;
        RECT 131.215 212.415 131.615 213.215 ;
        RECT 131.785 213.945 132.740 214.165 ;
        RECT 133.055 214.015 133.720 214.190 ;
        RECT 133.925 214.015 134.255 214.795 ;
        RECT 131.785 213.045 131.995 213.945 ;
        RECT 132.165 213.215 132.855 213.775 ;
        RECT 131.785 212.875 132.740 213.045 ;
        RECT 132.015 212.245 132.285 212.705 ;
        RECT 132.455 212.415 132.740 212.875 ;
        RECT 133.055 212.985 133.395 214.015 ;
        RECT 134.425 213.825 134.695 214.595 ;
        RECT 133.565 213.655 134.695 213.825 ;
        RECT 134.865 213.705 138.375 214.795 ;
        RECT 138.545 213.705 139.755 214.795 ;
        RECT 140.040 214.165 140.325 214.625 ;
        RECT 140.495 214.335 140.765 214.795 ;
        RECT 140.040 213.945 140.995 214.165 ;
        RECT 133.565 213.155 133.815 213.655 ;
        RECT 133.055 212.815 133.740 212.985 ;
        RECT 133.995 212.905 134.355 213.485 ;
        RECT 133.030 212.245 133.365 212.645 ;
        RECT 133.535 212.415 133.740 212.815 ;
        RECT 134.525 212.745 134.695 213.655 ;
        RECT 133.950 212.245 134.225 212.725 ;
        RECT 134.435 212.415 134.695 212.745 ;
        RECT 134.865 213.015 136.515 213.535 ;
        RECT 136.685 213.185 138.375 213.705 ;
        RECT 134.865 212.245 138.375 213.015 ;
        RECT 138.545 212.995 139.065 213.535 ;
        RECT 139.235 213.165 139.755 213.705 ;
        RECT 139.925 213.215 140.615 213.775 ;
        RECT 140.785 213.045 140.995 213.945 ;
        RECT 138.545 212.245 139.755 212.995 ;
        RECT 140.040 212.875 140.995 213.045 ;
        RECT 141.165 213.775 141.565 214.625 ;
        RECT 141.755 214.165 142.035 214.625 ;
        RECT 142.555 214.335 142.880 214.795 ;
        RECT 141.755 213.945 142.880 214.165 ;
        RECT 141.165 213.215 142.260 213.775 ;
        RECT 142.430 213.485 142.880 213.945 ;
        RECT 143.050 213.655 143.435 214.625 ;
        RECT 140.040 212.415 140.325 212.875 ;
        RECT 140.495 212.245 140.765 212.705 ;
        RECT 141.165 212.415 141.565 213.215 ;
        RECT 142.430 213.155 142.985 213.485 ;
        RECT 142.430 213.045 142.880 213.155 ;
        RECT 141.755 212.875 142.880 213.045 ;
        RECT 143.155 212.985 143.435 213.655 ;
        RECT 144.525 213.630 144.815 214.795 ;
        RECT 145.075 213.865 145.245 214.625 ;
        RECT 145.425 214.035 145.755 214.795 ;
        RECT 145.075 213.695 145.740 213.865 ;
        RECT 145.925 213.720 146.195 214.625 ;
        RECT 145.570 213.550 145.740 213.695 ;
        RECT 145.005 213.145 145.335 213.515 ;
        RECT 145.570 213.220 145.855 213.550 ;
        RECT 141.755 212.415 142.035 212.875 ;
        RECT 142.555 212.245 142.880 212.705 ;
        RECT 143.050 212.415 143.435 212.985 ;
        RECT 144.525 212.245 144.815 212.970 ;
        RECT 145.570 212.965 145.740 213.220 ;
        RECT 145.075 212.795 145.740 212.965 ;
        RECT 146.025 212.920 146.195 213.720 ;
        RECT 145.075 212.415 145.245 212.795 ;
        RECT 145.425 212.245 145.755 212.625 ;
        RECT 145.935 212.415 146.195 212.920 ;
        RECT 146.365 213.720 146.635 214.625 ;
        RECT 146.805 214.035 147.135 214.795 ;
        RECT 147.315 213.865 147.485 214.625 ;
        RECT 146.365 212.920 146.535 213.720 ;
        RECT 146.820 213.695 147.485 213.865 ;
        RECT 147.745 213.705 151.255 214.795 ;
        RECT 146.820 213.550 146.990 213.695 ;
        RECT 146.705 213.220 146.990 213.550 ;
        RECT 146.820 212.965 146.990 213.220 ;
        RECT 147.225 213.145 147.555 213.515 ;
        RECT 147.745 213.015 149.395 213.535 ;
        RECT 149.565 213.185 151.255 213.705 ;
        RECT 152.345 213.720 152.615 214.625 ;
        RECT 152.785 214.035 153.115 214.795 ;
        RECT 153.295 213.865 153.465 214.625 ;
        RECT 146.365 212.415 146.625 212.920 ;
        RECT 146.820 212.795 147.485 212.965 ;
        RECT 146.805 212.245 147.135 212.625 ;
        RECT 147.315 212.415 147.485 212.795 ;
        RECT 147.745 212.245 151.255 213.015 ;
        RECT 152.345 212.920 152.515 213.720 ;
        RECT 152.800 213.695 153.465 213.865 ;
        RECT 153.725 213.705 156.315 214.795 ;
        RECT 152.800 213.550 152.970 213.695 ;
        RECT 152.685 213.220 152.970 213.550 ;
        RECT 152.800 212.965 152.970 213.220 ;
        RECT 153.205 213.145 153.535 213.515 ;
        RECT 153.725 213.015 154.935 213.535 ;
        RECT 155.105 213.185 156.315 213.705 ;
        RECT 156.945 213.705 158.155 214.795 ;
        RECT 156.945 213.165 157.465 213.705 ;
        RECT 152.345 212.415 152.605 212.920 ;
        RECT 152.800 212.795 153.465 212.965 ;
        RECT 152.785 212.245 153.115 212.625 ;
        RECT 153.295 212.415 153.465 212.795 ;
        RECT 153.725 212.245 156.315 213.015 ;
        RECT 157.635 212.995 158.155 213.535 ;
        RECT 156.945 212.245 158.155 212.995 ;
        RECT 2.760 212.075 158.240 212.245 ;
        RECT 2.845 211.325 4.055 212.075 ;
        RECT 2.845 210.785 3.365 211.325 ;
        RECT 4.225 211.305 7.735 212.075 ;
        RECT 7.905 211.325 9.115 212.075 ;
        RECT 9.335 211.420 9.665 211.855 ;
        RECT 9.835 211.465 10.005 212.075 ;
        RECT 9.285 211.335 9.665 211.420 ;
        RECT 10.175 211.335 10.505 211.860 ;
        RECT 10.765 211.545 10.975 212.075 ;
        RECT 11.250 211.625 12.035 211.795 ;
        RECT 12.205 211.625 12.610 211.795 ;
        RECT 3.535 210.615 4.055 211.155 ;
        RECT 4.225 210.785 5.875 211.305 ;
        RECT 6.045 210.615 7.735 211.135 ;
        RECT 7.905 210.785 8.425 211.325 ;
        RECT 9.285 211.295 9.510 211.335 ;
        RECT 8.595 210.615 9.115 211.155 ;
        RECT 2.845 209.525 4.055 210.615 ;
        RECT 4.225 209.525 7.735 210.615 ;
        RECT 7.905 209.525 9.115 210.615 ;
        RECT 9.285 210.715 9.455 211.295 ;
        RECT 10.175 211.165 10.375 211.335 ;
        RECT 11.250 211.165 11.420 211.625 ;
        RECT 9.625 210.835 10.375 211.165 ;
        RECT 10.545 210.835 11.420 211.165 ;
        RECT 9.285 210.665 9.500 210.715 ;
        RECT 9.285 210.585 9.675 210.665 ;
        RECT 9.345 209.740 9.675 210.585 ;
        RECT 10.185 210.630 10.375 210.835 ;
        RECT 9.845 209.525 10.015 210.535 ;
        RECT 10.185 210.255 11.080 210.630 ;
        RECT 10.185 209.695 10.525 210.255 ;
        RECT 10.755 209.525 11.070 210.025 ;
        RECT 11.250 209.995 11.420 210.835 ;
        RECT 11.590 211.125 12.055 211.455 ;
        RECT 12.440 211.395 12.610 211.625 ;
        RECT 12.790 211.575 13.160 212.075 ;
        RECT 13.480 211.625 14.155 211.795 ;
        RECT 14.350 211.625 14.685 211.795 ;
        RECT 11.590 210.165 11.910 211.125 ;
        RECT 12.440 211.095 13.270 211.395 ;
        RECT 12.080 210.195 12.270 210.915 ;
        RECT 12.440 210.025 12.610 211.095 ;
        RECT 13.070 211.065 13.270 211.095 ;
        RECT 12.780 210.845 12.950 210.915 ;
        RECT 13.480 210.845 13.650 211.625 ;
        RECT 14.515 211.485 14.685 211.625 ;
        RECT 14.855 211.615 15.105 212.075 ;
        RECT 12.780 210.675 13.650 210.845 ;
        RECT 13.820 211.205 14.345 211.425 ;
        RECT 14.515 211.355 14.740 211.485 ;
        RECT 12.780 210.585 13.290 210.675 ;
        RECT 11.250 209.825 12.135 209.995 ;
        RECT 12.360 209.695 12.610 210.025 ;
        RECT 12.780 209.525 12.950 210.325 ;
        RECT 13.120 209.970 13.290 210.585 ;
        RECT 13.820 210.505 13.990 211.205 ;
        RECT 13.460 210.140 13.990 210.505 ;
        RECT 14.160 210.440 14.400 211.035 ;
        RECT 14.570 210.250 14.740 211.355 ;
        RECT 14.910 210.495 15.190 211.445 ;
        RECT 14.435 210.120 14.740 210.250 ;
        RECT 13.120 209.800 14.225 209.970 ;
        RECT 14.435 209.695 14.685 210.120 ;
        RECT 14.855 209.525 15.120 209.985 ;
        RECT 15.360 209.695 15.545 211.815 ;
        RECT 15.715 211.695 16.045 212.075 ;
        RECT 16.215 211.525 16.385 211.815 ;
        RECT 15.720 211.355 16.385 211.525 ;
        RECT 17.220 211.445 17.505 211.905 ;
        RECT 17.675 211.615 17.945 212.075 ;
        RECT 15.720 210.365 15.950 211.355 ;
        RECT 17.220 211.275 18.175 211.445 ;
        RECT 16.120 210.535 16.470 211.185 ;
        RECT 17.105 210.545 17.795 211.105 ;
        RECT 17.965 210.375 18.175 211.275 ;
        RECT 15.720 210.195 16.385 210.365 ;
        RECT 15.715 209.525 16.045 210.025 ;
        RECT 16.215 209.695 16.385 210.195 ;
        RECT 17.220 210.155 18.175 210.375 ;
        RECT 18.345 211.105 18.745 211.905 ;
        RECT 18.935 211.445 19.215 211.905 ;
        RECT 19.735 211.615 20.060 212.075 ;
        RECT 18.935 211.275 20.060 211.445 ;
        RECT 20.230 211.335 20.615 211.905 ;
        RECT 20.785 211.530 26.130 212.075 ;
        RECT 19.610 211.165 20.060 211.275 ;
        RECT 18.345 210.545 19.440 211.105 ;
        RECT 19.610 210.835 20.165 211.165 ;
        RECT 17.220 209.695 17.505 210.155 ;
        RECT 17.675 209.525 17.945 209.985 ;
        RECT 18.345 209.695 18.745 210.545 ;
        RECT 19.610 210.375 20.060 210.835 ;
        RECT 20.335 210.665 20.615 211.335 ;
        RECT 22.370 210.700 22.710 211.530 ;
        RECT 26.305 211.305 27.975 212.075 ;
        RECT 28.605 211.350 28.895 212.075 ;
        RECT 29.065 211.530 34.410 212.075 ;
        RECT 34.585 211.530 39.930 212.075 ;
        RECT 40.105 211.530 45.450 212.075 ;
        RECT 45.625 211.530 50.970 212.075 ;
        RECT 18.935 210.155 20.060 210.375 ;
        RECT 18.935 209.695 19.215 210.155 ;
        RECT 19.735 209.525 20.060 209.985 ;
        RECT 20.230 209.695 20.615 210.665 ;
        RECT 24.190 209.960 24.540 211.210 ;
        RECT 26.305 210.785 27.055 211.305 ;
        RECT 27.225 210.615 27.975 211.135 ;
        RECT 30.650 210.700 30.990 211.530 ;
        RECT 20.785 209.525 26.130 209.960 ;
        RECT 26.305 209.525 27.975 210.615 ;
        RECT 28.605 209.525 28.895 210.690 ;
        RECT 32.470 209.960 32.820 211.210 ;
        RECT 36.170 210.700 36.510 211.530 ;
        RECT 37.990 209.960 38.340 211.210 ;
        RECT 41.690 210.700 42.030 211.530 ;
        RECT 43.510 209.960 43.860 211.210 ;
        RECT 47.210 210.700 47.550 211.530 ;
        RECT 51.145 211.305 53.735 212.075 ;
        RECT 54.365 211.350 54.655 212.075 ;
        RECT 54.825 211.305 56.495 212.075 ;
        RECT 49.030 209.960 49.380 211.210 ;
        RECT 51.145 210.785 52.355 211.305 ;
        RECT 52.525 210.615 53.735 211.135 ;
        RECT 54.825 210.785 55.575 211.305 ;
        RECT 57.125 211.255 57.385 212.075 ;
        RECT 57.555 211.255 57.885 211.675 ;
        RECT 58.065 211.590 58.855 211.855 ;
        RECT 57.635 211.165 57.885 211.255 ;
        RECT 29.065 209.525 34.410 209.960 ;
        RECT 34.585 209.525 39.930 209.960 ;
        RECT 40.105 209.525 45.450 209.960 ;
        RECT 45.625 209.525 50.970 209.960 ;
        RECT 51.145 209.525 53.735 210.615 ;
        RECT 54.365 209.525 54.655 210.690 ;
        RECT 55.745 210.615 56.495 211.135 ;
        RECT 54.825 209.525 56.495 210.615 ;
        RECT 57.125 210.205 57.465 211.085 ;
        RECT 57.635 210.915 58.430 211.165 ;
        RECT 57.125 209.525 57.385 210.035 ;
        RECT 57.635 209.695 57.805 210.915 ;
        RECT 58.600 210.735 58.855 211.590 ;
        RECT 59.025 211.435 59.225 211.855 ;
        RECT 59.415 211.615 59.745 212.075 ;
        RECT 59.025 210.915 59.435 211.435 ;
        RECT 59.915 211.425 60.175 211.905 ;
        RECT 59.605 210.735 59.835 211.165 ;
        RECT 58.045 210.565 59.835 210.735 ;
        RECT 58.045 210.200 58.295 210.565 ;
        RECT 58.465 210.205 58.795 210.395 ;
        RECT 59.015 210.270 59.730 210.565 ;
        RECT 60.005 210.395 60.175 211.425 ;
        RECT 58.465 210.030 58.660 210.205 ;
        RECT 58.045 209.525 58.660 210.030 ;
        RECT 58.830 209.695 59.305 210.035 ;
        RECT 59.475 209.525 59.690 210.070 ;
        RECT 59.900 209.695 60.175 210.395 ;
        RECT 60.345 209.695 60.605 211.905 ;
        RECT 60.775 211.695 61.105 212.075 ;
        RECT 61.315 211.165 61.510 211.740 ;
        RECT 61.780 211.165 61.965 211.745 ;
        RECT 60.775 210.245 60.945 211.165 ;
        RECT 61.255 210.835 61.510 211.165 ;
        RECT 61.735 210.835 61.965 211.165 ;
        RECT 62.215 211.735 63.695 211.905 ;
        RECT 62.215 210.835 62.385 211.735 ;
        RECT 62.555 211.235 63.105 211.565 ;
        RECT 63.295 211.405 63.695 211.735 ;
        RECT 63.875 211.695 64.205 212.075 ;
        RECT 64.515 211.575 64.775 211.905 ;
        RECT 61.315 210.525 61.510 210.835 ;
        RECT 61.780 210.525 61.965 210.835 ;
        RECT 62.555 210.245 62.725 211.235 ;
        RECT 63.295 210.925 63.465 211.405 ;
        RECT 64.045 211.215 64.255 211.395 ;
        RECT 63.635 211.045 64.255 211.215 ;
        RECT 60.775 210.075 62.725 210.245 ;
        RECT 62.895 210.755 63.465 210.925 ;
        RECT 64.605 210.875 64.775 211.575 ;
        RECT 64.945 211.425 65.205 211.870 ;
        RECT 65.480 211.595 65.650 212.075 ;
        RECT 65.860 211.425 66.190 211.875 ;
        RECT 66.360 211.595 66.530 212.075 ;
        RECT 66.715 211.575 66.950 211.905 ;
        RECT 67.120 211.675 67.450 212.075 ;
        RECT 66.715 211.425 66.885 211.575 ;
        RECT 67.620 211.505 67.790 211.855 ;
        RECT 67.960 211.675 68.350 212.075 ;
        RECT 68.520 211.555 68.775 211.855 ;
        RECT 68.520 211.505 68.915 211.555 ;
        RECT 67.110 211.440 68.915 211.505 ;
        RECT 64.945 211.255 65.625 211.425 ;
        RECT 62.895 210.245 63.065 210.755 ;
        RECT 63.645 210.705 64.775 210.875 ;
        RECT 63.645 210.585 63.815 210.705 ;
        RECT 63.235 210.415 63.815 210.585 ;
        RECT 62.895 210.075 63.635 210.245 ;
        RECT 64.085 210.205 64.435 210.535 ;
        RECT 60.775 209.525 61.105 209.905 ;
        RECT 61.530 209.695 61.700 210.075 ;
        RECT 61.960 209.525 62.290 209.905 ;
        RECT 62.485 209.695 62.655 210.075 ;
        RECT 62.865 209.525 63.195 209.905 ;
        RECT 63.445 209.695 63.635 210.075 ;
        RECT 64.605 210.025 64.775 210.705 ;
        RECT 64.945 210.520 65.285 211.085 ;
        RECT 65.455 210.350 65.625 211.255 ;
        RECT 65.795 211.255 66.885 211.425 ;
        RECT 67.055 211.335 68.915 211.440 ;
        RECT 67.055 211.270 67.260 211.335 ;
        RECT 65.795 210.745 65.965 211.255 ;
        RECT 67.055 211.085 67.225 211.270 ;
        RECT 66.135 210.915 67.225 211.085 ;
        RECT 67.395 210.745 67.580 211.165 ;
        RECT 65.795 210.460 67.080 210.745 ;
        RECT 67.260 210.460 67.580 210.745 ;
        RECT 67.750 210.460 68.060 211.165 ;
        RECT 68.250 210.835 68.540 211.165 ;
        RECT 63.875 209.525 64.205 209.905 ;
        RECT 64.515 209.695 64.775 210.025 ;
        RECT 64.945 210.290 65.625 210.350 ;
        RECT 68.250 210.290 68.480 210.835 ;
        RECT 64.945 210.120 68.480 210.290 ;
        RECT 64.945 209.940 65.205 210.120 ;
        RECT 68.710 209.950 68.915 211.335 ;
        RECT 69.085 211.325 70.295 212.075 ;
        RECT 70.465 211.575 70.805 212.075 ;
        RECT 69.085 210.785 69.605 211.325 ;
        RECT 69.775 210.615 70.295 211.155 ;
        RECT 70.465 210.835 70.805 211.405 ;
        RECT 70.975 211.165 71.220 211.855 ;
        RECT 71.415 211.575 71.745 212.075 ;
        RECT 71.945 211.505 72.115 211.855 ;
        RECT 72.290 211.675 72.620 212.075 ;
        RECT 72.790 211.505 72.960 211.855 ;
        RECT 73.130 211.675 73.510 212.075 ;
        RECT 71.945 211.335 73.530 211.505 ;
        RECT 73.700 211.400 73.975 211.745 ;
        RECT 73.360 211.165 73.530 211.335 ;
        RECT 70.975 210.835 71.630 211.165 ;
        RECT 70.525 210.795 70.695 210.835 ;
        RECT 65.410 209.525 65.770 209.950 ;
        RECT 66.280 209.525 66.610 209.950 ;
        RECT 67.115 209.525 67.455 209.950 ;
        RECT 68.380 209.735 68.915 209.950 ;
        RECT 69.085 209.525 70.295 210.615 ;
        RECT 70.465 209.525 70.805 210.600 ;
        RECT 70.975 210.240 71.215 210.835 ;
        RECT 71.410 210.375 71.730 210.665 ;
        RECT 71.900 210.545 72.640 211.165 ;
        RECT 72.810 210.835 73.190 211.165 ;
        RECT 73.360 210.835 73.635 211.165 ;
        RECT 73.360 210.665 73.530 210.835 ;
        RECT 73.805 210.665 73.975 211.400 ;
        RECT 74.145 211.305 75.815 212.075 ;
        RECT 74.145 210.785 74.895 211.305 ;
        RECT 75.990 211.255 76.265 212.075 ;
        RECT 76.435 211.435 76.765 211.905 ;
        RECT 76.935 211.605 77.105 212.075 ;
        RECT 77.275 211.435 77.605 211.905 ;
        RECT 77.775 211.605 77.945 212.075 ;
        RECT 78.115 211.435 78.445 211.905 ;
        RECT 78.615 211.605 78.785 212.075 ;
        RECT 78.955 211.435 79.285 211.905 ;
        RECT 79.455 211.605 79.740 212.075 ;
        RECT 76.435 211.255 79.955 211.435 ;
        RECT 80.125 211.350 80.415 212.075 ;
        RECT 80.585 211.615 81.145 211.905 ;
        RECT 81.315 211.615 81.565 212.075 ;
        RECT 72.870 210.495 73.530 210.665 ;
        RECT 72.870 210.375 73.040 210.495 ;
        RECT 71.410 210.205 73.040 210.375 ;
        RECT 70.990 209.745 73.040 210.035 ;
        RECT 73.210 209.525 73.490 210.325 ;
        RECT 73.700 209.695 73.975 210.665 ;
        RECT 75.065 210.615 75.815 211.135 ;
        RECT 76.040 210.885 77.700 211.085 ;
        RECT 78.020 210.885 79.385 211.085 ;
        RECT 79.555 210.715 79.955 211.255 ;
        RECT 74.145 209.525 75.815 210.615 ;
        RECT 75.990 210.495 78.025 210.705 ;
        RECT 75.990 209.695 76.265 210.495 ;
        RECT 76.435 209.525 76.765 210.325 ;
        RECT 76.935 209.695 77.105 210.495 ;
        RECT 77.275 209.525 77.525 210.325 ;
        RECT 77.695 209.865 78.025 210.495 ;
        RECT 78.195 210.415 79.955 210.715 ;
        RECT 78.195 210.035 78.365 210.415 ;
        RECT 78.535 209.865 78.865 210.225 ;
        RECT 79.035 210.035 79.205 210.415 ;
        RECT 79.375 209.865 79.790 210.245 ;
        RECT 77.695 209.695 79.790 209.865 ;
        RECT 80.125 209.525 80.415 210.690 ;
        RECT 80.585 210.245 80.835 211.615 ;
        RECT 82.185 211.445 82.515 211.805 ;
        RECT 83.125 211.605 83.295 212.075 ;
        RECT 81.125 211.255 82.515 211.445 ;
        RECT 83.465 211.425 83.795 211.895 ;
        RECT 83.965 211.605 84.135 212.075 ;
        RECT 84.305 211.425 84.635 211.895 ;
        RECT 84.805 211.605 85.505 212.075 ;
        RECT 85.675 211.435 86.005 211.905 ;
        RECT 86.175 211.605 86.345 212.075 ;
        RECT 86.515 211.435 86.855 211.905 ;
        RECT 87.025 211.530 92.370 212.075 ;
        RECT 82.885 211.255 84.635 211.425 ;
        RECT 84.850 211.255 86.855 211.435 ;
        RECT 81.125 211.165 81.295 211.255 ;
        RECT 81.005 210.835 81.295 211.165 ;
        RECT 81.465 210.835 81.805 211.085 ;
        RECT 82.025 210.835 82.700 211.085 ;
        RECT 81.125 210.585 81.295 210.835 ;
        RECT 81.565 210.795 81.735 210.835 ;
        RECT 81.125 210.415 82.065 210.585 ;
        RECT 82.435 210.475 82.700 210.835 ;
        RECT 82.885 210.705 83.175 211.255 ;
        RECT 84.850 211.085 85.070 211.255 ;
        RECT 83.345 210.915 85.070 211.085 ;
        RECT 82.885 210.535 84.595 210.705 ;
        RECT 82.485 210.455 82.655 210.475 ;
        RECT 80.585 209.695 81.045 210.245 ;
        RECT 81.235 209.525 81.565 210.245 ;
        RECT 81.765 209.865 82.065 210.415 ;
        RECT 82.235 209.525 82.515 210.195 ;
        RECT 83.085 209.525 83.335 210.365 ;
        RECT 83.505 209.695 83.755 210.535 ;
        RECT 84.325 210.455 84.595 210.535 ;
        RECT 84.850 210.665 85.070 210.915 ;
        RECT 85.240 210.835 85.715 211.085 ;
        RECT 85.885 210.835 86.345 211.085 ;
        RECT 86.515 210.835 86.855 211.085 ;
        RECT 84.850 210.495 85.940 210.665 ;
        RECT 83.925 209.525 84.175 210.365 ;
        RECT 84.345 209.695 84.595 210.455 ;
        RECT 84.805 209.525 85.505 210.325 ;
        RECT 85.675 209.865 85.940 210.495 ;
        RECT 86.110 210.110 86.345 210.835 ;
        RECT 88.610 210.700 88.950 211.530 ;
        RECT 92.545 211.305 96.055 212.075 ;
        RECT 97.345 211.445 97.675 211.805 ;
        RECT 98.295 211.615 98.545 212.075 ;
        RECT 98.715 211.615 99.275 211.905 ;
        RECT 86.515 209.865 86.855 210.665 ;
        RECT 90.430 209.960 90.780 211.210 ;
        RECT 92.545 210.785 94.195 211.305 ;
        RECT 97.345 211.255 98.735 211.445 ;
        RECT 98.565 211.165 98.735 211.255 ;
        RECT 94.365 210.615 96.055 211.135 ;
        RECT 85.675 209.695 86.855 209.865 ;
        RECT 87.025 209.525 92.370 209.960 ;
        RECT 92.545 209.525 96.055 210.615 ;
        RECT 97.160 210.835 97.835 211.085 ;
        RECT 98.055 210.835 98.395 211.085 ;
        RECT 98.565 210.835 98.855 211.165 ;
        RECT 97.160 210.475 97.425 210.835 ;
        RECT 98.125 210.795 98.295 210.835 ;
        RECT 98.565 210.585 98.735 210.835 ;
        RECT 97.205 210.455 97.375 210.475 ;
        RECT 97.795 210.415 98.735 210.585 ;
        RECT 97.345 209.525 97.625 210.195 ;
        RECT 97.795 209.865 98.095 210.415 ;
        RECT 99.025 210.245 99.275 211.615 ;
        RECT 98.295 209.525 98.625 210.245 ;
        RECT 98.815 209.695 99.275 210.245 ;
        RECT 99.445 211.400 99.705 211.905 ;
        RECT 99.885 211.695 100.215 212.075 ;
        RECT 100.395 211.525 100.565 211.905 ;
        RECT 99.445 210.600 99.615 211.400 ;
        RECT 99.900 211.355 100.565 211.525 ;
        RECT 100.825 211.575 101.085 211.905 ;
        RECT 101.295 211.595 101.570 212.075 ;
        RECT 99.900 211.100 100.070 211.355 ;
        RECT 99.785 210.770 100.070 211.100 ;
        RECT 100.305 210.805 100.635 211.175 ;
        RECT 99.900 210.625 100.070 210.770 ;
        RECT 100.825 210.665 100.995 211.575 ;
        RECT 101.780 211.505 101.985 211.905 ;
        RECT 102.155 211.675 102.490 212.075 ;
        RECT 101.165 210.835 101.525 211.415 ;
        RECT 101.780 211.335 102.465 211.505 ;
        RECT 101.705 210.665 101.955 211.165 ;
        RECT 99.445 209.695 99.715 210.600 ;
        RECT 99.900 210.455 100.565 210.625 ;
        RECT 99.885 209.525 100.215 210.285 ;
        RECT 100.395 209.695 100.565 210.455 ;
        RECT 100.825 210.495 101.955 210.665 ;
        RECT 100.825 209.725 101.095 210.495 ;
        RECT 102.125 210.305 102.465 211.335 ;
        RECT 102.865 211.445 103.195 211.805 ;
        RECT 103.815 211.615 104.065 212.075 ;
        RECT 104.235 211.615 104.795 211.905 ;
        RECT 102.865 211.255 104.255 211.445 ;
        RECT 104.085 211.165 104.255 211.255 ;
        RECT 102.680 210.835 103.355 211.085 ;
        RECT 103.575 210.835 103.915 211.085 ;
        RECT 104.085 210.835 104.375 211.165 ;
        RECT 102.680 210.475 102.945 210.835 ;
        RECT 103.185 210.795 103.355 210.835 ;
        RECT 103.645 210.795 103.815 210.835 ;
        RECT 104.085 210.585 104.255 210.835 ;
        RECT 101.265 209.525 101.595 210.305 ;
        RECT 101.800 210.130 102.465 210.305 ;
        RECT 103.315 210.415 104.255 210.585 ;
        RECT 101.800 209.725 101.985 210.130 ;
        RECT 102.155 209.525 102.490 209.950 ;
        RECT 102.865 209.525 103.145 210.195 ;
        RECT 103.315 209.865 103.615 210.415 ;
        RECT 104.545 210.245 104.795 211.615 ;
        RECT 105.885 211.350 106.175 212.075 ;
        RECT 103.815 209.525 104.145 210.245 ;
        RECT 104.335 209.695 104.795 210.245 ;
        RECT 105.885 209.525 106.175 210.690 ;
        RECT 106.355 209.705 106.615 211.895 ;
        RECT 106.875 211.705 107.545 212.075 ;
        RECT 107.725 211.525 108.035 211.895 ;
        RECT 106.805 211.325 108.035 211.525 ;
        RECT 106.805 210.655 107.095 211.325 ;
        RECT 108.215 211.145 108.445 211.785 ;
        RECT 108.625 211.345 108.915 212.075 ;
        RECT 109.105 211.415 109.380 212.075 ;
        RECT 109.550 211.445 109.800 211.905 ;
        RECT 109.975 211.580 110.305 212.075 ;
        RECT 109.550 211.235 109.720 211.445 ;
        RECT 110.485 211.410 110.715 211.855 ;
        RECT 107.275 210.835 107.740 211.145 ;
        RECT 107.920 210.835 108.445 211.145 ;
        RECT 108.625 210.835 108.925 211.165 ;
        RECT 109.105 210.715 109.720 211.235 ;
        RECT 109.890 210.735 110.120 211.165 ;
        RECT 110.305 210.915 110.715 211.410 ;
        RECT 110.885 211.590 111.675 211.855 ;
        RECT 110.885 210.735 111.140 211.590 ;
        RECT 111.310 210.915 111.695 211.395 ;
        RECT 111.875 211.265 112.145 212.075 ;
        RECT 112.315 211.265 112.645 211.905 ;
        RECT 112.815 211.265 113.055 212.075 ;
        RECT 111.865 210.835 112.215 211.085 ;
        RECT 106.805 210.435 107.575 210.655 ;
        RECT 106.785 209.525 107.125 210.255 ;
        RECT 107.305 209.705 107.575 210.435 ;
        RECT 107.755 210.415 108.915 210.655 ;
        RECT 107.755 209.705 107.985 210.415 ;
        RECT 108.155 209.525 108.485 210.235 ;
        RECT 108.655 209.705 108.915 210.415 ;
        RECT 109.105 209.525 109.365 210.535 ;
        RECT 109.535 210.365 109.705 210.715 ;
        RECT 109.890 210.565 111.680 210.735 ;
        RECT 112.385 210.665 112.555 211.265 ;
        RECT 112.725 210.835 113.075 211.085 ;
        RECT 109.535 209.695 109.810 210.365 ;
        RECT 110.010 209.525 110.225 210.370 ;
        RECT 110.450 210.270 110.700 210.565 ;
        RECT 110.925 210.205 111.255 210.395 ;
        RECT 110.410 209.695 110.885 210.035 ;
        RECT 111.065 210.030 111.255 210.205 ;
        RECT 111.425 210.200 111.680 210.565 ;
        RECT 111.065 209.525 111.695 210.030 ;
        RECT 111.875 209.525 112.205 210.665 ;
        RECT 112.385 210.495 113.065 210.665 ;
        RECT 113.725 210.495 113.955 211.835 ;
        RECT 114.135 210.995 114.365 211.895 ;
        RECT 114.565 211.295 114.810 212.075 ;
        RECT 114.980 211.535 115.410 211.895 ;
        RECT 115.990 211.705 116.720 212.075 ;
        RECT 114.980 211.345 116.720 211.535 ;
        RECT 114.980 211.115 115.200 211.345 ;
        RECT 112.735 209.710 113.065 210.495 ;
        RECT 114.135 210.315 114.475 210.995 ;
        RECT 113.725 210.115 114.475 210.315 ;
        RECT 114.655 210.815 115.200 211.115 ;
        RECT 113.725 209.725 113.965 210.115 ;
        RECT 114.135 209.525 114.485 209.935 ;
        RECT 114.655 209.705 114.985 210.815 ;
        RECT 115.370 210.545 115.795 211.165 ;
        RECT 115.990 210.545 116.250 211.165 ;
        RECT 116.460 210.835 116.720 211.345 ;
        RECT 115.155 210.175 116.180 210.375 ;
        RECT 115.155 209.705 115.335 210.175 ;
        RECT 115.505 209.525 115.835 210.005 ;
        RECT 116.010 209.705 116.180 210.175 ;
        RECT 116.445 209.525 116.730 210.665 ;
        RECT 116.920 209.705 117.200 211.895 ;
        RECT 117.385 211.305 120.895 212.075 ;
        RECT 121.065 211.325 122.275 212.075 ;
        RECT 122.535 211.525 122.705 211.815 ;
        RECT 122.875 211.695 123.205 212.075 ;
        RECT 122.535 211.355 123.200 211.525 ;
        RECT 117.385 210.785 119.035 211.305 ;
        RECT 119.205 210.615 120.895 211.135 ;
        RECT 121.065 210.785 121.585 211.325 ;
        RECT 121.755 210.615 122.275 211.155 ;
        RECT 117.385 209.525 120.895 210.615 ;
        RECT 121.065 209.525 122.275 210.615 ;
        RECT 122.450 210.535 122.800 211.185 ;
        RECT 122.970 210.365 123.200 211.355 ;
        RECT 122.535 210.195 123.200 210.365 ;
        RECT 122.535 209.695 122.705 210.195 ;
        RECT 122.875 209.525 123.205 210.025 ;
        RECT 123.375 209.695 123.560 211.815 ;
        RECT 123.815 211.615 124.065 212.075 ;
        RECT 124.235 211.625 124.570 211.795 ;
        RECT 124.765 211.625 125.440 211.795 ;
        RECT 124.235 211.485 124.405 211.625 ;
        RECT 123.730 210.495 124.010 211.445 ;
        RECT 124.180 211.355 124.405 211.485 ;
        RECT 124.180 210.250 124.350 211.355 ;
        RECT 124.575 211.205 125.100 211.425 ;
        RECT 124.520 210.440 124.760 211.035 ;
        RECT 124.930 210.505 125.100 211.205 ;
        RECT 125.270 210.845 125.440 211.625 ;
        RECT 125.760 211.575 126.130 212.075 ;
        RECT 126.310 211.625 126.715 211.795 ;
        RECT 126.885 211.625 127.670 211.795 ;
        RECT 126.310 211.395 126.480 211.625 ;
        RECT 125.650 211.095 126.480 211.395 ;
        RECT 126.865 211.125 127.330 211.455 ;
        RECT 125.650 211.065 125.850 211.095 ;
        RECT 125.970 210.845 126.140 210.915 ;
        RECT 125.270 210.675 126.140 210.845 ;
        RECT 125.630 210.585 126.140 210.675 ;
        RECT 124.180 210.120 124.485 210.250 ;
        RECT 124.930 210.140 125.460 210.505 ;
        RECT 123.800 209.525 124.065 209.985 ;
        RECT 124.235 209.695 124.485 210.120 ;
        RECT 125.630 209.970 125.800 210.585 ;
        RECT 124.695 209.800 125.800 209.970 ;
        RECT 125.970 209.525 126.140 210.325 ;
        RECT 126.310 210.025 126.480 211.095 ;
        RECT 126.650 210.195 126.840 210.915 ;
        RECT 127.010 210.165 127.330 211.125 ;
        RECT 127.500 211.165 127.670 211.625 ;
        RECT 127.945 211.545 128.155 212.075 ;
        RECT 128.415 211.335 128.745 211.860 ;
        RECT 128.915 211.465 129.085 212.075 ;
        RECT 129.255 211.420 129.585 211.855 ;
        RECT 129.255 211.335 129.635 211.420 ;
        RECT 128.545 211.165 128.745 211.335 ;
        RECT 129.410 211.295 129.635 211.335 ;
        RECT 127.500 210.835 128.375 211.165 ;
        RECT 128.545 210.835 129.295 211.165 ;
        RECT 126.310 209.695 126.560 210.025 ;
        RECT 127.500 209.995 127.670 210.835 ;
        RECT 128.545 210.630 128.735 210.835 ;
        RECT 129.465 210.715 129.635 211.295 ;
        RECT 129.805 211.305 131.475 212.075 ;
        RECT 131.645 211.350 131.935 212.075 ;
        RECT 132.105 211.335 132.490 211.905 ;
        RECT 132.660 211.615 132.985 212.075 ;
        RECT 133.505 211.445 133.785 211.905 ;
        RECT 129.805 210.785 130.555 211.305 ;
        RECT 129.420 210.665 129.635 210.715 ;
        RECT 127.840 210.255 128.735 210.630 ;
        RECT 129.245 210.585 129.635 210.665 ;
        RECT 130.725 210.615 131.475 211.135 ;
        RECT 126.785 209.825 127.670 209.995 ;
        RECT 127.850 209.525 128.165 210.025 ;
        RECT 128.395 209.695 128.735 210.255 ;
        RECT 128.905 209.525 129.075 210.535 ;
        RECT 129.245 209.740 129.575 210.585 ;
        RECT 129.805 209.525 131.475 210.615 ;
        RECT 131.645 209.525 131.935 210.690 ;
        RECT 132.105 210.665 132.385 211.335 ;
        RECT 132.660 211.275 133.785 211.445 ;
        RECT 132.660 211.165 133.110 211.275 ;
        RECT 132.555 210.835 133.110 211.165 ;
        RECT 133.975 211.105 134.375 211.905 ;
        RECT 134.775 211.615 135.045 212.075 ;
        RECT 135.215 211.445 135.500 211.905 ;
        RECT 135.785 211.530 141.130 212.075 ;
        RECT 141.305 211.530 146.650 212.075 ;
        RECT 146.825 211.530 152.170 212.075 ;
        RECT 132.105 209.695 132.490 210.665 ;
        RECT 132.660 210.375 133.110 210.835 ;
        RECT 133.280 210.545 134.375 211.105 ;
        RECT 132.660 210.155 133.785 210.375 ;
        RECT 132.660 209.525 132.985 209.985 ;
        RECT 133.505 209.695 133.785 210.155 ;
        RECT 133.975 209.695 134.375 210.545 ;
        RECT 134.545 211.275 135.500 211.445 ;
        RECT 134.545 210.375 134.755 211.275 ;
        RECT 134.925 210.545 135.615 211.105 ;
        RECT 137.370 210.700 137.710 211.530 ;
        RECT 134.545 210.155 135.500 210.375 ;
        RECT 134.775 209.525 135.045 209.985 ;
        RECT 135.215 209.695 135.500 210.155 ;
        RECT 139.190 209.960 139.540 211.210 ;
        RECT 142.890 210.700 143.230 211.530 ;
        RECT 144.710 209.960 145.060 211.210 ;
        RECT 148.410 210.700 148.750 211.530 ;
        RECT 152.345 211.305 155.855 212.075 ;
        RECT 156.945 211.325 158.155 212.075 ;
        RECT 150.230 209.960 150.580 211.210 ;
        RECT 152.345 210.785 153.995 211.305 ;
        RECT 154.165 210.615 155.855 211.135 ;
        RECT 135.785 209.525 141.130 209.960 ;
        RECT 141.305 209.525 146.650 209.960 ;
        RECT 146.825 209.525 152.170 209.960 ;
        RECT 152.345 209.525 155.855 210.615 ;
        RECT 156.945 210.615 157.465 211.155 ;
        RECT 157.635 210.785 158.155 211.325 ;
        RECT 156.945 209.525 158.155 210.615 ;
        RECT 2.760 209.355 158.240 209.525 ;
        RECT 2.845 208.265 4.055 209.355 ;
        RECT 4.225 208.920 9.570 209.355 ;
        RECT 2.845 207.555 3.365 208.095 ;
        RECT 3.535 207.725 4.055 208.265 ;
        RECT 2.845 206.805 4.055 207.555 ;
        RECT 5.810 207.350 6.150 208.180 ;
        RECT 7.630 207.670 7.980 208.920 ;
        RECT 10.665 207.635 11.185 209.185 ;
        RECT 11.355 208.630 11.685 209.355 ;
        RECT 12.160 208.725 12.445 209.185 ;
        RECT 12.615 208.895 12.885 209.355 ;
        RECT 12.160 208.505 13.115 208.725 ;
        RECT 4.225 206.805 9.570 207.350 ;
        RECT 10.845 206.805 11.185 207.465 ;
        RECT 11.355 206.975 11.875 208.460 ;
        RECT 12.045 207.775 12.735 208.335 ;
        RECT 12.905 207.605 13.115 208.505 ;
        RECT 12.160 207.435 13.115 207.605 ;
        RECT 13.285 208.335 13.685 209.185 ;
        RECT 13.875 208.725 14.155 209.185 ;
        RECT 14.675 208.895 15.000 209.355 ;
        RECT 13.875 208.505 15.000 208.725 ;
        RECT 13.285 207.775 14.380 208.335 ;
        RECT 14.550 208.045 15.000 208.505 ;
        RECT 15.170 208.215 15.555 209.185 ;
        RECT 12.160 206.975 12.445 207.435 ;
        RECT 12.615 206.805 12.885 207.265 ;
        RECT 13.285 206.975 13.685 207.775 ;
        RECT 14.550 207.715 15.105 208.045 ;
        RECT 14.550 207.605 15.000 207.715 ;
        RECT 13.875 207.435 15.000 207.605 ;
        RECT 15.275 207.545 15.555 208.215 ;
        RECT 15.725 208.190 16.015 209.355 ;
        RECT 16.185 208.265 18.775 209.355 ;
        RECT 19.495 208.685 19.665 209.185 ;
        RECT 19.835 208.855 20.165 209.355 ;
        RECT 19.495 208.515 20.160 208.685 ;
        RECT 13.875 206.975 14.155 207.435 ;
        RECT 14.675 206.805 15.000 207.265 ;
        RECT 15.170 206.975 15.555 207.545 ;
        RECT 16.185 207.575 17.395 208.095 ;
        RECT 17.565 207.745 18.775 208.265 ;
        RECT 19.410 207.695 19.760 208.345 ;
        RECT 15.725 206.805 16.015 207.530 ;
        RECT 16.185 206.805 18.775 207.575 ;
        RECT 19.930 207.525 20.160 208.515 ;
        RECT 19.495 207.355 20.160 207.525 ;
        RECT 19.495 207.065 19.665 207.355 ;
        RECT 19.835 206.805 20.165 207.185 ;
        RECT 20.335 207.065 20.520 209.185 ;
        RECT 20.760 208.895 21.025 209.355 ;
        RECT 21.195 208.760 21.445 209.185 ;
        RECT 21.655 208.910 22.760 209.080 ;
        RECT 21.140 208.630 21.445 208.760 ;
        RECT 20.690 207.435 20.970 208.385 ;
        RECT 21.140 207.525 21.310 208.630 ;
        RECT 21.480 207.845 21.720 208.440 ;
        RECT 21.890 208.375 22.420 208.740 ;
        RECT 21.890 207.675 22.060 208.375 ;
        RECT 22.590 208.295 22.760 208.910 ;
        RECT 22.930 208.555 23.100 209.355 ;
        RECT 23.270 208.855 23.520 209.185 ;
        RECT 23.745 208.885 24.630 209.055 ;
        RECT 22.590 208.205 23.100 208.295 ;
        RECT 21.140 207.395 21.365 207.525 ;
        RECT 21.535 207.455 22.060 207.675 ;
        RECT 22.230 208.035 23.100 208.205 ;
        RECT 20.775 206.805 21.025 207.265 ;
        RECT 21.195 207.255 21.365 207.395 ;
        RECT 22.230 207.255 22.400 208.035 ;
        RECT 22.930 207.965 23.100 208.035 ;
        RECT 22.610 207.785 22.810 207.815 ;
        RECT 23.270 207.785 23.440 208.855 ;
        RECT 23.610 207.965 23.800 208.685 ;
        RECT 22.610 207.485 23.440 207.785 ;
        RECT 23.970 207.755 24.290 208.715 ;
        RECT 21.195 207.085 21.530 207.255 ;
        RECT 21.725 207.085 22.400 207.255 ;
        RECT 22.720 206.805 23.090 207.305 ;
        RECT 23.270 207.255 23.440 207.485 ;
        RECT 23.825 207.425 24.290 207.755 ;
        RECT 24.460 208.045 24.630 208.885 ;
        RECT 24.810 208.855 25.125 209.355 ;
        RECT 25.355 208.625 25.695 209.185 ;
        RECT 24.800 208.250 25.695 208.625 ;
        RECT 25.865 208.345 26.035 209.355 ;
        RECT 25.505 208.045 25.695 208.250 ;
        RECT 26.205 208.295 26.535 209.140 ;
        RECT 26.705 208.440 26.875 209.355 ;
        RECT 26.205 208.215 26.595 208.295 ;
        RECT 27.225 208.265 29.815 209.355 ;
        RECT 30.100 208.725 30.385 209.185 ;
        RECT 30.555 208.895 30.825 209.355 ;
        RECT 30.100 208.505 31.055 208.725 ;
        RECT 26.380 208.165 26.595 208.215 ;
        RECT 24.460 207.715 25.335 208.045 ;
        RECT 25.505 207.715 26.255 208.045 ;
        RECT 24.460 207.255 24.630 207.715 ;
        RECT 25.505 207.545 25.705 207.715 ;
        RECT 26.425 207.585 26.595 208.165 ;
        RECT 26.370 207.565 26.595 207.585 ;
        RECT 26.365 207.545 26.595 207.565 ;
        RECT 23.270 207.085 23.675 207.255 ;
        RECT 23.845 207.085 24.630 207.255 ;
        RECT 24.905 206.805 25.115 207.335 ;
        RECT 25.375 207.020 25.705 207.545 ;
        RECT 26.215 207.460 26.595 207.545 ;
        RECT 27.225 207.575 28.435 208.095 ;
        RECT 28.605 207.745 29.815 208.265 ;
        RECT 29.985 207.775 30.675 208.335 ;
        RECT 30.845 207.605 31.055 208.505 ;
        RECT 25.875 206.805 26.045 207.415 ;
        RECT 26.215 207.025 26.545 207.460 ;
        RECT 26.715 206.805 26.885 207.320 ;
        RECT 27.225 206.805 29.815 207.575 ;
        RECT 30.100 207.435 31.055 207.605 ;
        RECT 31.225 208.335 31.625 209.185 ;
        RECT 31.815 208.725 32.095 209.185 ;
        RECT 32.615 208.895 32.940 209.355 ;
        RECT 31.815 208.505 32.940 208.725 ;
        RECT 31.225 207.775 32.320 208.335 ;
        RECT 32.490 208.045 32.940 208.505 ;
        RECT 33.110 208.215 33.495 209.185 ;
        RECT 33.665 208.920 39.010 209.355 ;
        RECT 30.100 206.975 30.385 207.435 ;
        RECT 30.555 206.805 30.825 207.265 ;
        RECT 31.225 206.975 31.625 207.775 ;
        RECT 32.490 207.715 33.045 208.045 ;
        RECT 32.490 207.605 32.940 207.715 ;
        RECT 31.815 207.435 32.940 207.605 ;
        RECT 33.215 207.545 33.495 208.215 ;
        RECT 31.815 206.975 32.095 207.435 ;
        RECT 32.615 206.805 32.940 207.265 ;
        RECT 33.110 206.975 33.495 207.545 ;
        RECT 35.250 207.350 35.590 208.180 ;
        RECT 37.070 207.670 37.420 208.920 ;
        RECT 39.185 208.265 40.855 209.355 ;
        RECT 39.185 207.575 39.935 208.095 ;
        RECT 40.105 207.745 40.855 208.265 ;
        RECT 41.485 208.190 41.775 209.355 ;
        RECT 41.945 208.920 47.290 209.355 ;
        RECT 47.465 208.920 52.810 209.355 ;
        RECT 52.985 208.920 58.330 209.355 ;
        RECT 58.670 209.015 60.765 209.185 ;
        RECT 33.665 206.805 39.010 207.350 ;
        RECT 39.185 206.805 40.855 207.575 ;
        RECT 41.485 206.805 41.775 207.530 ;
        RECT 43.530 207.350 43.870 208.180 ;
        RECT 45.350 207.670 45.700 208.920 ;
        RECT 49.050 207.350 49.390 208.180 ;
        RECT 50.870 207.670 51.220 208.920 ;
        RECT 54.570 207.350 54.910 208.180 ;
        RECT 56.390 207.670 56.740 208.920 ;
        RECT 58.670 208.635 59.085 209.015 ;
        RECT 59.255 208.465 59.425 208.845 ;
        RECT 59.595 208.655 59.925 209.015 ;
        RECT 60.095 208.465 60.265 208.845 ;
        RECT 58.505 208.165 60.265 208.465 ;
        RECT 60.435 208.385 60.765 209.015 ;
        RECT 60.935 208.555 61.185 209.355 ;
        RECT 61.355 208.385 61.525 209.185 ;
        RECT 61.695 208.555 62.025 209.355 ;
        RECT 62.195 208.385 62.470 209.185 ;
        RECT 62.810 209.015 64.905 209.185 ;
        RECT 62.810 208.635 63.225 209.015 ;
        RECT 63.395 208.465 63.565 208.845 ;
        RECT 63.735 208.655 64.065 209.015 ;
        RECT 64.235 208.465 64.405 208.845 ;
        RECT 60.435 208.175 62.470 208.385 ;
        RECT 62.645 208.165 64.405 208.465 ;
        RECT 64.575 208.385 64.905 209.015 ;
        RECT 65.075 208.555 65.325 209.355 ;
        RECT 65.495 208.385 65.665 209.185 ;
        RECT 65.835 208.555 66.165 209.355 ;
        RECT 66.335 208.385 66.610 209.185 ;
        RECT 64.575 208.175 66.610 208.385 ;
        RECT 67.245 208.190 67.535 209.355 ;
        RECT 67.765 208.215 67.975 209.355 ;
        RECT 68.145 208.205 68.475 209.185 ;
        RECT 68.645 208.215 68.875 209.355 ;
        RECT 69.550 208.215 69.905 209.355 ;
        RECT 70.095 208.385 70.425 209.185 ;
        RECT 70.595 208.555 70.765 209.355 ;
        RECT 70.935 208.385 71.265 209.185 ;
        RECT 71.435 208.555 71.605 209.355 ;
        RECT 71.775 208.385 72.105 209.185 ;
        RECT 72.275 208.555 72.445 209.355 ;
        RECT 72.615 208.385 72.945 209.185 ;
        RECT 73.115 208.555 73.285 209.355 ;
        RECT 73.455 208.385 73.785 209.185 ;
        RECT 73.955 208.555 74.125 209.355 ;
        RECT 74.295 208.385 74.625 209.185 ;
        RECT 74.795 208.555 74.965 209.355 ;
        RECT 75.135 208.385 75.465 209.185 ;
        RECT 75.635 208.555 75.805 209.355 ;
        RECT 75.975 208.385 76.305 209.185 ;
        RECT 58.505 207.625 58.905 208.165 ;
        RECT 59.075 207.795 60.440 207.995 ;
        RECT 60.760 207.795 62.420 207.995 ;
        RECT 62.645 207.625 63.045 208.165 ;
        RECT 63.215 207.795 64.580 207.995 ;
        RECT 64.900 207.795 66.560 207.995 ;
        RECT 58.505 207.445 62.025 207.625 ;
        RECT 41.945 206.805 47.290 207.350 ;
        RECT 47.465 206.805 52.810 207.350 ;
        RECT 52.985 206.805 58.330 207.350 ;
        RECT 58.720 206.805 59.005 207.275 ;
        RECT 59.175 206.975 59.505 207.445 ;
        RECT 59.675 206.805 59.845 207.275 ;
        RECT 60.015 206.975 60.345 207.445 ;
        RECT 60.515 206.805 60.685 207.275 ;
        RECT 60.855 206.975 61.185 207.445 ;
        RECT 61.355 206.805 61.525 207.275 ;
        RECT 61.695 206.975 62.025 207.445 ;
        RECT 62.195 206.805 62.470 207.625 ;
        RECT 62.645 207.445 66.165 207.625 ;
        RECT 62.860 206.805 63.145 207.275 ;
        RECT 63.315 206.975 63.645 207.445 ;
        RECT 63.815 206.805 63.985 207.275 ;
        RECT 64.155 206.975 64.485 207.445 ;
        RECT 64.655 206.805 64.825 207.275 ;
        RECT 64.995 206.975 65.325 207.445 ;
        RECT 65.495 206.805 65.665 207.275 ;
        RECT 65.835 206.975 66.165 207.445 ;
        RECT 66.335 206.805 66.610 207.625 ;
        RECT 67.245 206.805 67.535 207.530 ;
        RECT 67.765 206.805 67.975 207.625 ;
        RECT 68.145 207.605 68.395 208.205 ;
        RECT 70.095 208.185 76.305 208.385 ;
        RECT 76.475 208.215 76.730 209.355 ;
        RECT 77.105 208.685 77.385 209.355 ;
        RECT 77.555 208.465 77.855 209.015 ;
        RECT 78.055 208.635 78.385 209.355 ;
        RECT 78.575 208.635 79.035 209.185 ;
        RECT 68.565 207.795 68.895 208.045 ;
        RECT 70.095 207.625 70.345 208.185 ;
        RECT 70.515 207.795 72.530 207.995 ;
        RECT 72.700 207.795 73.180 208.185 ;
        RECT 76.920 208.045 77.185 208.405 ;
        RECT 77.555 208.295 78.495 208.465 ;
        RECT 78.325 208.045 78.495 208.295 ;
        RECT 73.455 207.795 76.310 208.015 ;
        RECT 76.920 207.795 77.595 208.045 ;
        RECT 77.815 207.795 78.155 208.045 ;
        RECT 72.700 207.625 72.945 207.795 ;
        RECT 78.325 207.715 78.615 208.045 ;
        RECT 78.325 207.625 78.495 207.715 ;
        RECT 68.145 206.975 68.475 207.605 ;
        RECT 68.645 206.805 68.875 207.625 ;
        RECT 69.550 207.205 69.925 207.625 ;
        RECT 70.095 207.375 72.945 207.625 ;
        RECT 73.115 207.455 76.730 207.625 ;
        RECT 73.115 207.205 73.365 207.455 ;
        RECT 69.550 206.975 73.365 207.205 ;
        RECT 73.535 206.805 73.705 207.285 ;
        RECT 73.875 206.975 74.205 207.455 ;
        RECT 74.375 206.805 74.545 207.285 ;
        RECT 74.715 206.975 75.045 207.455 ;
        RECT 75.215 206.805 75.385 207.285 ;
        RECT 75.555 206.975 75.885 207.455 ;
        RECT 76.055 206.805 76.225 207.285 ;
        RECT 76.395 206.975 76.730 207.455 ;
        RECT 77.105 207.435 78.495 207.625 ;
        RECT 77.105 207.075 77.435 207.435 ;
        RECT 78.785 207.265 79.035 208.635 ;
        RECT 79.205 208.265 80.415 209.355 ;
        RECT 78.055 206.805 78.305 207.265 ;
        RECT 78.475 206.975 79.035 207.265 ;
        RECT 79.205 207.555 79.725 208.095 ;
        RECT 79.895 207.725 80.415 208.265 ;
        RECT 80.585 208.930 81.120 209.145 ;
        RECT 82.045 208.930 82.385 209.355 ;
        RECT 82.890 208.930 83.220 209.355 ;
        RECT 83.730 208.930 84.090 209.355 ;
        RECT 79.205 206.805 80.415 207.555 ;
        RECT 80.585 207.545 80.790 208.930 ;
        RECT 84.295 208.760 84.555 208.940 ;
        RECT 81.020 208.590 84.555 208.760 ;
        RECT 84.925 208.685 85.205 209.355 ;
        RECT 81.020 208.045 81.250 208.590 ;
        RECT 83.875 208.530 84.555 208.590 ;
        RECT 80.960 207.715 81.250 208.045 ;
        RECT 81.440 207.715 81.750 208.420 ;
        RECT 81.920 208.135 82.240 208.420 ;
        RECT 82.420 208.135 83.705 208.420 ;
        RECT 81.920 207.715 82.105 208.135 ;
        RECT 82.275 207.795 83.365 207.965 ;
        RECT 82.275 207.610 82.445 207.795 ;
        RECT 83.535 207.625 83.705 208.135 ;
        RECT 82.240 207.545 82.445 207.610 ;
        RECT 80.585 207.440 82.445 207.545 ;
        RECT 82.615 207.455 83.705 207.625 ;
        RECT 83.875 207.625 84.045 208.530 ;
        RECT 85.375 208.465 85.675 209.015 ;
        RECT 85.875 208.635 86.205 209.355 ;
        RECT 86.395 208.635 86.855 209.185 ;
        RECT 84.215 207.795 84.555 208.360 ;
        RECT 84.740 208.045 85.005 208.405 ;
        RECT 85.375 208.295 86.315 208.465 ;
        RECT 86.145 208.045 86.315 208.295 ;
        RECT 84.740 207.795 85.415 208.045 ;
        RECT 85.635 207.795 85.975 208.045 ;
        RECT 86.145 207.715 86.435 208.045 ;
        RECT 86.145 207.625 86.315 207.715 ;
        RECT 83.875 207.455 84.555 207.625 ;
        RECT 80.585 207.375 82.390 207.440 ;
        RECT 80.585 207.325 80.980 207.375 ;
        RECT 80.725 207.025 80.980 207.325 ;
        RECT 81.150 206.805 81.540 207.205 ;
        RECT 81.710 207.025 81.880 207.375 ;
        RECT 82.615 207.305 82.785 207.455 ;
        RECT 82.050 206.805 82.380 207.205 ;
        RECT 82.550 206.975 82.785 207.305 ;
        RECT 82.970 206.805 83.140 207.285 ;
        RECT 83.310 207.005 83.640 207.455 ;
        RECT 83.850 206.805 84.020 207.285 ;
        RECT 84.295 207.010 84.555 207.455 ;
        RECT 84.925 207.435 86.315 207.625 ;
        RECT 84.925 207.075 85.255 207.435 ;
        RECT 86.605 207.265 86.855 208.635 ;
        RECT 87.025 208.265 89.615 209.355 ;
        RECT 89.985 208.685 90.265 209.355 ;
        RECT 90.435 208.465 90.735 209.015 ;
        RECT 90.935 208.635 91.265 209.355 ;
        RECT 91.455 208.635 91.915 209.185 ;
        RECT 85.875 206.805 86.125 207.265 ;
        RECT 86.295 206.975 86.855 207.265 ;
        RECT 87.025 207.575 88.235 208.095 ;
        RECT 88.405 207.745 89.615 208.265 ;
        RECT 89.800 208.045 90.065 208.405 ;
        RECT 90.435 208.295 91.375 208.465 ;
        RECT 91.205 208.045 91.375 208.295 ;
        RECT 89.800 207.795 90.475 208.045 ;
        RECT 90.695 207.795 91.035 208.045 ;
        RECT 91.205 207.715 91.495 208.045 ;
        RECT 91.205 207.625 91.375 207.715 ;
        RECT 87.025 206.805 89.615 207.575 ;
        RECT 89.985 207.435 91.375 207.625 ;
        RECT 89.985 207.075 90.315 207.435 ;
        RECT 91.665 207.265 91.915 208.635 ;
        RECT 93.005 208.190 93.295 209.355 ;
        RECT 93.465 208.265 96.055 209.355 ;
        RECT 96.425 208.685 96.705 209.355 ;
        RECT 96.875 208.465 97.175 209.015 ;
        RECT 97.375 208.635 97.705 209.355 ;
        RECT 97.895 208.635 98.355 209.185 ;
        RECT 93.465 207.575 94.675 208.095 ;
        RECT 94.845 207.745 96.055 208.265 ;
        RECT 96.240 208.045 96.505 208.405 ;
        RECT 96.875 208.295 97.815 208.465 ;
        RECT 97.205 208.045 97.375 208.075 ;
        RECT 97.645 208.045 97.815 208.295 ;
        RECT 96.240 207.795 96.915 208.045 ;
        RECT 97.135 207.795 97.475 208.045 ;
        RECT 97.645 207.715 97.935 208.045 ;
        RECT 97.645 207.625 97.815 207.715 ;
        RECT 90.935 206.805 91.185 207.265 ;
        RECT 91.355 206.975 91.915 207.265 ;
        RECT 93.005 206.805 93.295 207.530 ;
        RECT 93.465 206.805 96.055 207.575 ;
        RECT 96.425 207.435 97.815 207.625 ;
        RECT 96.425 207.075 96.755 207.435 ;
        RECT 98.105 207.265 98.355 208.635 ;
        RECT 98.530 208.685 98.785 209.185 ;
        RECT 98.955 208.855 99.285 209.355 ;
        RECT 98.530 208.515 99.280 208.685 ;
        RECT 98.530 207.695 98.880 208.345 ;
        RECT 99.050 207.525 99.280 208.515 ;
        RECT 97.375 206.805 97.625 207.265 ;
        RECT 97.795 206.975 98.355 207.265 ;
        RECT 98.530 207.355 99.280 207.525 ;
        RECT 98.530 207.065 98.785 207.355 ;
        RECT 98.955 206.805 99.285 207.185 ;
        RECT 99.455 207.065 99.625 209.185 ;
        RECT 99.795 208.385 100.120 209.170 ;
        RECT 100.290 208.895 100.540 209.355 ;
        RECT 100.710 208.855 100.960 209.185 ;
        RECT 101.175 208.855 101.855 209.185 ;
        RECT 100.710 208.725 100.880 208.855 ;
        RECT 100.485 208.555 100.880 208.725 ;
        RECT 99.855 207.335 100.315 208.385 ;
        RECT 100.485 207.195 100.655 208.555 ;
        RECT 101.050 208.295 101.515 208.685 ;
        RECT 100.825 207.485 101.175 208.105 ;
        RECT 101.345 207.705 101.515 208.295 ;
        RECT 101.685 208.075 101.855 208.855 ;
        RECT 102.025 208.755 102.195 209.095 ;
        RECT 102.430 208.925 102.760 209.355 ;
        RECT 102.930 208.755 103.100 209.095 ;
        RECT 103.395 208.895 103.765 209.355 ;
        RECT 102.025 208.585 103.100 208.755 ;
        RECT 103.935 208.725 104.105 209.185 ;
        RECT 104.340 208.845 105.210 209.185 ;
        RECT 105.380 208.895 105.630 209.355 ;
        RECT 103.545 208.555 104.105 208.725 ;
        RECT 103.545 208.415 103.715 208.555 ;
        RECT 102.215 208.245 103.715 208.415 ;
        RECT 104.410 208.385 104.870 208.675 ;
        RECT 101.685 207.905 103.375 208.075 ;
        RECT 101.345 207.485 101.700 207.705 ;
        RECT 101.870 207.195 102.040 207.905 ;
        RECT 102.245 207.485 103.035 207.735 ;
        RECT 103.205 207.725 103.375 207.905 ;
        RECT 103.545 207.555 103.715 208.245 ;
        RECT 99.985 206.805 100.315 207.165 ;
        RECT 100.485 207.025 100.980 207.195 ;
        RECT 101.185 207.025 102.040 207.195 ;
        RECT 102.915 206.805 103.245 207.265 ;
        RECT 103.455 207.165 103.715 207.555 ;
        RECT 103.905 208.375 104.870 208.385 ;
        RECT 105.040 208.465 105.210 208.845 ;
        RECT 105.800 208.805 105.970 209.095 ;
        RECT 106.150 208.975 106.480 209.355 ;
        RECT 105.800 208.635 106.600 208.805 ;
        RECT 103.905 208.215 104.580 208.375 ;
        RECT 105.040 208.295 106.260 208.465 ;
        RECT 103.905 207.425 104.115 208.215 ;
        RECT 105.040 208.205 105.210 208.295 ;
        RECT 104.285 207.425 104.635 208.045 ;
        RECT 104.805 208.035 105.210 208.205 ;
        RECT 104.805 207.255 104.975 208.035 ;
        RECT 105.145 207.585 105.365 207.865 ;
        RECT 105.545 207.755 106.085 208.125 ;
        RECT 106.430 208.015 106.600 208.635 ;
        RECT 106.775 208.295 106.945 209.355 ;
        RECT 107.155 208.345 107.445 209.185 ;
        RECT 107.615 208.515 107.785 209.355 ;
        RECT 107.995 208.345 108.245 209.185 ;
        RECT 108.455 208.515 108.625 209.355 ;
        RECT 109.105 208.635 109.565 209.185 ;
        RECT 109.755 208.635 110.085 209.355 ;
        RECT 107.155 208.175 108.880 208.345 ;
        RECT 105.145 207.415 105.675 207.585 ;
        RECT 103.455 206.995 103.805 207.165 ;
        RECT 104.025 206.975 104.975 207.255 ;
        RECT 105.145 206.805 105.335 207.245 ;
        RECT 105.505 207.185 105.675 207.415 ;
        RECT 105.845 207.355 106.085 207.755 ;
        RECT 106.255 208.005 106.600 208.015 ;
        RECT 106.255 207.795 108.285 208.005 ;
        RECT 106.255 207.540 106.580 207.795 ;
        RECT 108.470 207.625 108.880 208.175 ;
        RECT 106.255 207.185 106.575 207.540 ;
        RECT 105.505 207.015 106.575 207.185 ;
        RECT 106.775 206.805 106.945 207.615 ;
        RECT 107.115 207.455 108.880 207.625 ;
        RECT 107.115 206.975 107.445 207.455 ;
        RECT 107.615 206.805 107.785 207.275 ;
        RECT 107.955 206.975 108.285 207.455 ;
        RECT 108.455 206.805 108.625 207.275 ;
        RECT 109.105 207.265 109.355 208.635 ;
        RECT 110.285 208.465 110.585 209.015 ;
        RECT 110.755 208.685 111.035 209.355 ;
        RECT 111.445 209.015 112.585 209.185 ;
        RECT 111.445 208.555 111.745 209.015 ;
        RECT 109.645 208.295 110.585 208.465 ;
        RECT 109.645 208.045 109.815 208.295 ;
        RECT 110.070 208.045 110.240 208.075 ;
        RECT 110.955 208.045 111.220 208.405 ;
        RECT 111.915 208.385 112.245 208.845 ;
        RECT 109.525 207.715 109.815 208.045 ;
        RECT 109.985 207.795 110.325 208.045 ;
        RECT 110.545 207.795 111.220 208.045 ;
        RECT 111.485 208.165 112.245 208.385 ;
        RECT 112.415 208.385 112.585 209.015 ;
        RECT 112.755 208.555 113.085 209.355 ;
        RECT 113.255 208.385 113.530 209.185 ;
        RECT 112.415 208.175 113.530 208.385 ;
        RECT 113.705 208.265 117.215 209.355 ;
        RECT 117.385 208.265 118.595 209.355 ;
        RECT 109.645 207.625 109.815 207.715 ;
        RECT 111.485 207.625 111.700 208.165 ;
        RECT 111.870 207.795 112.640 207.995 ;
        RECT 112.810 207.795 113.530 207.995 ;
        RECT 109.645 207.435 111.035 207.625 ;
        RECT 111.485 207.455 113.085 207.625 ;
        RECT 109.105 206.975 109.665 207.265 ;
        RECT 109.835 206.805 110.085 207.265 ;
        RECT 110.705 207.075 111.035 207.435 ;
        RECT 111.915 207.445 113.085 207.455 ;
        RECT 111.455 206.805 111.745 207.275 ;
        RECT 111.915 206.975 112.245 207.445 ;
        RECT 112.415 206.805 112.585 207.275 ;
        RECT 112.755 206.975 113.085 207.445 ;
        RECT 113.255 206.805 113.530 207.625 ;
        RECT 113.705 207.575 115.355 208.095 ;
        RECT 115.525 207.745 117.215 208.265 ;
        RECT 113.705 206.805 117.215 207.575 ;
        RECT 117.385 207.555 117.905 208.095 ;
        RECT 118.075 207.725 118.595 208.265 ;
        RECT 118.765 208.190 119.055 209.355 ;
        RECT 119.225 208.920 124.570 209.355 ;
        RECT 117.385 206.805 118.595 207.555 ;
        RECT 118.765 206.805 119.055 207.530 ;
        RECT 120.810 207.350 121.150 208.180 ;
        RECT 122.630 207.670 122.980 208.920 ;
        RECT 124.745 208.265 126.415 209.355 ;
        RECT 124.745 207.575 125.495 208.095 ;
        RECT 125.665 207.745 126.415 208.265 ;
        RECT 127.050 208.215 127.305 209.355 ;
        RECT 127.500 208.805 128.695 209.135 ;
        RECT 127.555 208.045 127.725 208.605 ;
        RECT 127.950 208.385 128.370 208.635 ;
        RECT 128.875 208.555 129.155 209.355 ;
        RECT 127.950 208.215 129.195 208.385 ;
        RECT 129.365 208.215 129.635 209.185 ;
        RECT 129.805 208.920 135.150 209.355 ;
        RECT 135.325 208.920 140.670 209.355 ;
        RECT 129.025 208.045 129.195 208.215 ;
        RECT 127.050 207.795 127.385 208.045 ;
        RECT 127.555 207.715 128.295 208.045 ;
        RECT 129.025 207.715 129.255 208.045 ;
        RECT 127.555 207.625 127.805 207.715 ;
        RECT 119.225 206.805 124.570 207.350 ;
        RECT 124.745 206.805 126.415 207.575 ;
        RECT 127.070 207.455 127.805 207.625 ;
        RECT 129.025 207.545 129.195 207.715 ;
        RECT 127.070 206.985 127.380 207.455 ;
        RECT 128.455 207.375 129.195 207.545 ;
        RECT 129.465 207.480 129.635 208.215 ;
        RECT 127.550 206.805 128.285 207.285 ;
        RECT 128.455 207.025 128.625 207.375 ;
        RECT 128.795 206.805 129.175 207.205 ;
        RECT 129.365 207.135 129.635 207.480 ;
        RECT 131.390 207.350 131.730 208.180 ;
        RECT 133.210 207.670 133.560 208.920 ;
        RECT 136.910 207.350 137.250 208.180 ;
        RECT 138.730 207.670 139.080 208.920 ;
        RECT 140.845 208.265 144.355 209.355 ;
        RECT 140.845 207.575 142.495 208.095 ;
        RECT 142.665 207.745 144.355 208.265 ;
        RECT 144.525 208.190 144.815 209.355 ;
        RECT 144.985 208.920 150.330 209.355 ;
        RECT 150.505 208.920 155.850 209.355 ;
        RECT 129.805 206.805 135.150 207.350 ;
        RECT 135.325 206.805 140.670 207.350 ;
        RECT 140.845 206.805 144.355 207.575 ;
        RECT 144.525 206.805 144.815 207.530 ;
        RECT 146.570 207.350 146.910 208.180 ;
        RECT 148.390 207.670 148.740 208.920 ;
        RECT 152.090 207.350 152.430 208.180 ;
        RECT 153.910 207.670 154.260 208.920 ;
        RECT 156.945 208.265 158.155 209.355 ;
        RECT 156.945 207.725 157.465 208.265 ;
        RECT 157.635 207.555 158.155 208.095 ;
        RECT 144.985 206.805 150.330 207.350 ;
        RECT 150.505 206.805 155.850 207.350 ;
        RECT 156.945 206.805 158.155 207.555 ;
        RECT 2.760 206.635 158.240 206.805 ;
        RECT 2.845 205.885 4.055 206.635 ;
        RECT 4.225 206.090 9.570 206.635 ;
        RECT 2.845 205.345 3.365 205.885 ;
        RECT 3.535 205.175 4.055 205.715 ;
        RECT 5.810 205.260 6.150 206.090 ;
        RECT 10.210 205.795 10.470 206.635 ;
        RECT 10.645 205.890 10.900 206.465 ;
        RECT 11.070 206.255 11.400 206.635 ;
        RECT 11.615 206.085 11.785 206.465 ;
        RECT 12.215 206.120 12.385 206.635 ;
        RECT 11.070 205.915 11.785 206.085 ;
        RECT 12.555 205.980 12.885 206.415 ;
        RECT 13.055 206.025 13.225 206.635 ;
        RECT 2.845 204.085 4.055 205.175 ;
        RECT 7.630 204.520 7.980 205.770 ;
        RECT 4.225 204.085 9.570 204.520 ;
        RECT 10.210 204.085 10.470 205.235 ;
        RECT 10.645 205.160 10.815 205.890 ;
        RECT 11.070 205.725 11.240 205.915 ;
        RECT 12.505 205.895 12.885 205.980 ;
        RECT 13.395 205.895 13.725 206.420 ;
        RECT 13.985 206.105 14.195 206.635 ;
        RECT 14.470 206.185 15.255 206.355 ;
        RECT 15.425 206.185 15.830 206.355 ;
        RECT 12.505 205.855 12.730 205.895 ;
        RECT 10.985 205.395 11.240 205.725 ;
        RECT 11.070 205.185 11.240 205.395 ;
        RECT 11.520 205.365 11.875 205.735 ;
        RECT 11.645 205.355 11.815 205.365 ;
        RECT 12.505 205.275 12.675 205.855 ;
        RECT 13.395 205.725 13.595 205.895 ;
        RECT 14.470 205.725 14.640 206.185 ;
        RECT 12.845 205.395 13.595 205.725 ;
        RECT 13.765 205.395 14.640 205.725 ;
        RECT 12.505 205.225 12.720 205.275 ;
        RECT 10.645 204.255 10.900 205.160 ;
        RECT 11.070 205.015 11.785 205.185 ;
        RECT 12.505 205.145 12.895 205.225 ;
        RECT 11.070 204.085 11.400 204.845 ;
        RECT 11.615 204.255 11.785 205.015 ;
        RECT 12.225 204.085 12.395 205.000 ;
        RECT 12.565 204.300 12.895 205.145 ;
        RECT 13.405 205.190 13.595 205.395 ;
        RECT 13.065 204.085 13.235 205.095 ;
        RECT 13.405 204.815 14.300 205.190 ;
        RECT 13.405 204.255 13.745 204.815 ;
        RECT 13.975 204.085 14.290 204.585 ;
        RECT 14.470 204.555 14.640 205.395 ;
        RECT 14.810 205.685 15.275 206.015 ;
        RECT 15.660 205.955 15.830 206.185 ;
        RECT 16.010 206.135 16.380 206.635 ;
        RECT 16.700 206.185 17.375 206.355 ;
        RECT 17.570 206.185 17.905 206.355 ;
        RECT 14.810 204.725 15.130 205.685 ;
        RECT 15.660 205.655 16.490 205.955 ;
        RECT 15.300 204.755 15.490 205.475 ;
        RECT 15.660 204.585 15.830 205.655 ;
        RECT 16.290 205.625 16.490 205.655 ;
        RECT 16.000 205.405 16.170 205.475 ;
        RECT 16.700 205.405 16.870 206.185 ;
        RECT 17.735 206.045 17.905 206.185 ;
        RECT 18.075 206.175 18.325 206.635 ;
        RECT 16.000 205.235 16.870 205.405 ;
        RECT 17.040 205.765 17.565 205.985 ;
        RECT 17.735 205.915 17.960 206.045 ;
        RECT 16.000 205.145 16.510 205.235 ;
        RECT 14.470 204.385 15.355 204.555 ;
        RECT 15.580 204.255 15.830 204.585 ;
        RECT 16.000 204.085 16.170 204.885 ;
        RECT 16.340 204.530 16.510 205.145 ;
        RECT 17.040 205.065 17.210 205.765 ;
        RECT 16.680 204.700 17.210 205.065 ;
        RECT 17.380 205.000 17.620 205.595 ;
        RECT 17.790 204.810 17.960 205.915 ;
        RECT 18.130 205.055 18.410 206.005 ;
        RECT 17.655 204.680 17.960 204.810 ;
        RECT 16.340 204.360 17.445 204.530 ;
        RECT 17.655 204.255 17.905 204.680 ;
        RECT 18.075 204.085 18.340 204.545 ;
        RECT 18.580 204.255 18.765 206.375 ;
        RECT 18.935 206.255 19.265 206.635 ;
        RECT 19.435 206.085 19.605 206.375 ;
        RECT 18.940 205.915 19.605 206.085 ;
        RECT 18.940 204.925 19.170 205.915 ;
        RECT 19.865 205.885 21.075 206.635 ;
        RECT 19.340 205.095 19.690 205.745 ;
        RECT 19.865 205.345 20.385 205.885 ;
        RECT 21.250 205.795 21.510 206.635 ;
        RECT 21.685 205.890 21.940 206.465 ;
        RECT 22.110 206.255 22.440 206.635 ;
        RECT 22.655 206.085 22.825 206.465 ;
        RECT 23.085 206.090 28.430 206.635 ;
        RECT 22.110 205.915 22.825 206.085 ;
        RECT 20.555 205.175 21.075 205.715 ;
        RECT 18.940 204.755 19.605 204.925 ;
        RECT 18.935 204.085 19.265 204.585 ;
        RECT 19.435 204.255 19.605 204.755 ;
        RECT 19.865 204.085 21.075 205.175 ;
        RECT 21.250 204.085 21.510 205.235 ;
        RECT 21.685 205.160 21.855 205.890 ;
        RECT 22.110 205.725 22.280 205.915 ;
        RECT 22.025 205.395 22.280 205.725 ;
        RECT 22.110 205.185 22.280 205.395 ;
        RECT 22.560 205.365 22.915 205.735 ;
        RECT 22.685 205.355 22.855 205.365 ;
        RECT 24.670 205.260 25.010 206.090 ;
        RECT 28.605 205.910 28.895 206.635 ;
        RECT 29.065 205.865 31.655 206.635 ;
        RECT 21.685 204.255 21.940 205.160 ;
        RECT 22.110 205.015 22.825 205.185 ;
        RECT 22.110 204.085 22.440 204.845 ;
        RECT 22.655 204.255 22.825 205.015 ;
        RECT 26.490 204.520 26.840 205.770 ;
        RECT 29.065 205.345 30.275 205.865 ;
        RECT 32.290 205.795 32.550 206.635 ;
        RECT 32.725 205.890 32.980 206.465 ;
        RECT 33.150 206.255 33.480 206.635 ;
        RECT 33.695 206.085 33.865 206.465 ;
        RECT 34.125 206.090 39.470 206.635 ;
        RECT 33.150 205.915 33.865 206.085 ;
        RECT 23.085 204.085 28.430 204.520 ;
        RECT 28.605 204.085 28.895 205.250 ;
        RECT 30.445 205.175 31.655 205.695 ;
        RECT 29.065 204.085 31.655 205.175 ;
        RECT 32.290 204.085 32.550 205.235 ;
        RECT 32.725 205.160 32.895 205.890 ;
        RECT 33.150 205.725 33.320 205.915 ;
        RECT 33.065 205.395 33.320 205.725 ;
        RECT 33.150 205.185 33.320 205.395 ;
        RECT 33.600 205.365 33.955 205.735 ;
        RECT 33.725 205.355 33.895 205.365 ;
        RECT 35.710 205.260 36.050 206.090 ;
        RECT 39.650 205.795 39.910 206.635 ;
        RECT 40.085 205.890 40.340 206.465 ;
        RECT 40.510 206.255 40.840 206.635 ;
        RECT 41.055 206.085 41.225 206.465 ;
        RECT 41.485 206.090 46.830 206.635 ;
        RECT 47.005 206.090 52.350 206.635 ;
        RECT 40.510 205.915 41.225 206.085 ;
        RECT 32.725 204.255 32.980 205.160 ;
        RECT 33.150 205.015 33.865 205.185 ;
        RECT 33.150 204.085 33.480 204.845 ;
        RECT 33.695 204.255 33.865 205.015 ;
        RECT 37.530 204.520 37.880 205.770 ;
        RECT 34.125 204.085 39.470 204.520 ;
        RECT 39.650 204.085 39.910 205.235 ;
        RECT 40.085 205.160 40.255 205.890 ;
        RECT 40.510 205.725 40.680 205.915 ;
        RECT 40.425 205.395 40.680 205.725 ;
        RECT 40.510 205.185 40.680 205.395 ;
        RECT 40.960 205.365 41.315 205.735 ;
        RECT 41.085 205.355 41.255 205.365 ;
        RECT 43.070 205.260 43.410 206.090 ;
        RECT 40.085 204.255 40.340 205.160 ;
        RECT 40.510 205.015 41.225 205.185 ;
        RECT 40.510 204.085 40.840 204.845 ;
        RECT 41.055 204.255 41.225 205.015 ;
        RECT 44.890 204.520 45.240 205.770 ;
        RECT 48.590 205.260 48.930 206.090 ;
        RECT 52.525 205.865 54.195 206.635 ;
        RECT 54.365 205.910 54.655 206.635 ;
        RECT 54.825 205.865 58.335 206.635 ;
        RECT 50.410 204.520 50.760 205.770 ;
        RECT 52.525 205.345 53.275 205.865 ;
        RECT 53.445 205.175 54.195 205.695 ;
        RECT 54.825 205.345 56.475 205.865 ;
        RECT 58.510 205.815 58.785 206.635 ;
        RECT 58.955 205.995 59.285 206.465 ;
        RECT 59.455 206.165 59.625 206.635 ;
        RECT 59.795 205.995 60.125 206.465 ;
        RECT 60.295 206.165 60.465 206.635 ;
        RECT 60.635 205.995 60.965 206.465 ;
        RECT 61.135 206.165 61.305 206.635 ;
        RECT 61.475 205.995 61.805 206.465 ;
        RECT 61.975 206.165 62.260 206.635 ;
        RECT 62.645 205.995 62.935 206.465 ;
        RECT 63.135 206.165 63.305 206.635 ;
        RECT 63.475 205.995 63.805 206.465 ;
        RECT 63.975 206.165 64.145 206.635 ;
        RECT 64.315 205.995 64.645 206.465 ;
        RECT 64.815 206.165 64.985 206.635 ;
        RECT 65.155 205.995 65.485 206.465 ;
        RECT 65.655 206.165 65.825 206.635 ;
        RECT 65.995 205.995 66.325 206.465 ;
        RECT 66.495 206.165 66.665 206.635 ;
        RECT 66.835 205.995 67.165 206.465 ;
        RECT 67.335 206.165 67.505 206.635 ;
        RECT 67.675 205.995 68.005 206.465 ;
        RECT 58.955 205.815 62.475 205.995 ;
        RECT 41.485 204.085 46.830 204.520 ;
        RECT 47.005 204.085 52.350 204.520 ;
        RECT 52.525 204.085 54.195 205.175 ;
        RECT 54.365 204.085 54.655 205.250 ;
        RECT 56.645 205.175 58.335 205.695 ;
        RECT 58.560 205.445 60.220 205.645 ;
        RECT 60.540 205.445 61.905 205.645 ;
        RECT 62.075 205.275 62.475 205.815 ;
        RECT 54.825 204.085 58.335 205.175 ;
        RECT 58.510 205.055 60.545 205.265 ;
        RECT 58.510 204.255 58.785 205.055 ;
        RECT 58.955 204.085 59.285 204.885 ;
        RECT 59.455 204.255 59.625 205.055 ;
        RECT 59.795 204.085 60.045 204.885 ;
        RECT 60.215 204.425 60.545 205.055 ;
        RECT 60.715 204.975 62.475 205.275 ;
        RECT 62.645 205.815 68.005 205.995 ;
        RECT 68.175 205.815 68.450 206.635 ;
        RECT 68.810 206.155 68.980 206.635 ;
        RECT 69.150 205.985 69.480 206.455 ;
        RECT 69.650 206.155 69.820 206.635 ;
        RECT 69.990 205.985 70.320 206.455 ;
        RECT 68.625 205.815 70.320 205.985 ;
        RECT 70.530 205.895 70.700 206.635 ;
        RECT 70.915 205.895 71.245 206.430 ;
        RECT 71.415 206.125 71.655 206.635 ;
        RECT 72.060 206.165 72.345 206.635 ;
        RECT 72.515 205.995 72.845 206.465 ;
        RECT 73.015 206.165 73.185 206.635 ;
        RECT 73.355 205.995 73.685 206.465 ;
        RECT 73.855 206.165 74.025 206.635 ;
        RECT 74.195 205.995 74.525 206.465 ;
        RECT 74.695 206.165 74.865 206.635 ;
        RECT 75.035 205.995 75.365 206.465 ;
        RECT 60.715 204.595 60.885 204.975 ;
        RECT 61.055 204.425 61.385 204.785 ;
        RECT 61.555 204.595 61.725 204.975 ;
        RECT 62.645 204.935 62.935 205.815 ;
        RECT 63.125 205.435 63.545 205.645 ;
        RECT 63.775 205.445 64.685 205.645 ;
        RECT 63.250 205.355 63.545 205.435 ;
        RECT 63.375 205.275 63.545 205.355 ;
        RECT 64.855 205.435 66.445 205.645 ;
        RECT 66.715 205.435 68.450 205.645 ;
        RECT 64.855 205.275 65.025 205.435 ;
        RECT 63.375 205.105 65.025 205.275 ;
        RECT 65.195 205.095 66.285 205.265 ;
        RECT 61.895 204.425 62.310 204.805 ;
        RECT 60.215 204.255 62.310 204.425 ;
        RECT 62.645 204.765 65.025 204.935 ;
        RECT 62.645 204.255 62.925 204.765 ;
        RECT 63.935 204.755 65.025 204.765 ;
        RECT 63.935 204.595 64.185 204.755 ;
        RECT 64.775 204.595 65.025 204.755 ;
        RECT 63.095 204.255 63.345 204.595 ;
        RECT 63.515 204.425 63.765 204.585 ;
        RECT 64.355 204.425 64.605 204.585 ;
        RECT 65.195 204.425 65.445 205.095 ;
        RECT 63.515 204.255 65.445 204.425 ;
        RECT 65.615 204.635 65.865 204.925 ;
        RECT 66.035 204.805 66.285 205.095 ;
        RECT 66.455 205.095 68.390 205.265 ;
        RECT 66.455 204.635 66.705 205.095 ;
        RECT 65.615 204.255 66.705 204.635 ;
        RECT 66.875 204.085 67.125 204.925 ;
        RECT 67.295 204.255 67.545 205.095 ;
        RECT 67.715 204.085 67.965 204.925 ;
        RECT 68.135 204.255 68.390 205.095 ;
        RECT 68.625 205.225 68.970 205.815 ;
        RECT 69.140 205.475 70.350 205.645 ;
        RECT 70.145 205.225 70.350 205.475 ;
        RECT 70.520 205.395 70.895 205.725 ;
        RECT 71.065 205.225 71.245 205.895 ;
        RECT 71.415 205.395 71.670 205.955 ;
        RECT 71.845 205.815 75.365 205.995 ;
        RECT 75.535 205.815 75.810 206.635 ;
        RECT 76.200 206.165 76.485 206.635 ;
        RECT 76.655 205.995 76.985 206.465 ;
        RECT 77.155 206.165 77.325 206.635 ;
        RECT 77.495 205.995 77.825 206.465 ;
        RECT 77.995 206.165 78.165 206.635 ;
        RECT 78.335 205.995 78.665 206.465 ;
        RECT 78.835 206.165 79.005 206.635 ;
        RECT 79.175 205.995 79.505 206.465 ;
        RECT 75.985 205.815 79.505 205.995 ;
        RECT 79.675 205.815 79.950 206.635 ;
        RECT 80.125 205.910 80.415 206.635 ;
        RECT 80.800 206.165 81.085 206.635 ;
        RECT 81.255 205.995 81.585 206.465 ;
        RECT 81.755 206.165 81.925 206.635 ;
        RECT 82.095 205.995 82.425 206.465 ;
        RECT 82.595 206.165 82.765 206.635 ;
        RECT 82.935 205.995 83.265 206.465 ;
        RECT 83.435 206.165 83.605 206.635 ;
        RECT 83.775 205.995 84.105 206.465 ;
        RECT 80.585 205.815 84.105 205.995 ;
        RECT 84.275 205.815 84.550 206.635 ;
        RECT 84.730 205.815 85.005 206.635 ;
        RECT 85.175 205.995 85.505 206.465 ;
        RECT 85.675 206.165 85.845 206.635 ;
        RECT 86.015 205.995 86.345 206.465 ;
        RECT 86.515 206.165 86.685 206.635 ;
        RECT 86.855 205.995 87.185 206.465 ;
        RECT 87.355 206.165 87.525 206.635 ;
        RECT 87.695 205.995 88.025 206.465 ;
        RECT 88.195 206.165 88.480 206.635 ;
        RECT 88.955 206.085 89.125 206.465 ;
        RECT 89.340 206.255 89.670 206.635 ;
        RECT 85.175 205.815 88.695 205.995 ;
        RECT 88.955 205.915 89.670 206.085 ;
        RECT 71.845 205.275 72.245 205.815 ;
        RECT 72.415 205.445 73.780 205.645 ;
        RECT 74.100 205.445 75.760 205.645 ;
        RECT 75.985 205.275 76.385 205.815 ;
        RECT 76.555 205.445 77.920 205.645 ;
        RECT 78.240 205.445 79.900 205.645 ;
        RECT 80.585 205.275 80.985 205.815 ;
        RECT 81.155 205.445 82.520 205.645 ;
        RECT 82.840 205.445 84.500 205.645 ;
        RECT 84.780 205.445 86.440 205.645 ;
        RECT 86.760 205.445 88.125 205.645 ;
        RECT 88.295 205.275 88.695 205.815 ;
        RECT 88.865 205.365 89.220 205.735 ;
        RECT 89.500 205.725 89.670 205.915 ;
        RECT 89.840 205.890 90.095 206.465 ;
        RECT 89.500 205.395 89.755 205.725 ;
        RECT 88.925 205.355 89.095 205.365 ;
        RECT 68.625 205.055 69.480 205.225 ;
        RECT 70.145 205.055 71.605 205.225 ;
        RECT 69.145 205.015 69.480 205.055 ;
        RECT 69.150 204.885 69.480 205.015 ;
        RECT 68.810 204.085 68.980 204.885 ;
        RECT 69.150 204.715 70.320 204.885 ;
        RECT 69.150 204.255 69.480 204.715 ;
        RECT 69.650 204.085 69.820 204.545 ;
        RECT 69.990 204.255 70.320 204.715 ;
        RECT 70.530 204.085 70.700 204.885 ;
        RECT 71.245 204.255 71.605 205.055 ;
        RECT 71.845 204.975 73.605 205.275 ;
        RECT 72.010 204.425 72.425 204.805 ;
        RECT 72.595 204.595 72.765 204.975 ;
        RECT 72.935 204.425 73.265 204.785 ;
        RECT 73.435 204.595 73.605 204.975 ;
        RECT 73.775 205.055 75.810 205.265 ;
        RECT 73.775 204.425 74.105 205.055 ;
        RECT 72.010 204.255 74.105 204.425 ;
        RECT 74.275 204.085 74.525 204.885 ;
        RECT 74.695 204.255 74.865 205.055 ;
        RECT 75.035 204.085 75.365 204.885 ;
        RECT 75.535 204.255 75.810 205.055 ;
        RECT 75.985 204.975 77.745 205.275 ;
        RECT 76.150 204.425 76.565 204.805 ;
        RECT 76.735 204.595 76.905 204.975 ;
        RECT 77.075 204.425 77.405 204.785 ;
        RECT 77.575 204.595 77.745 204.975 ;
        RECT 77.915 205.055 79.950 205.265 ;
        RECT 77.915 204.425 78.245 205.055 ;
        RECT 76.150 204.255 78.245 204.425 ;
        RECT 78.415 204.085 78.665 204.885 ;
        RECT 78.835 204.255 79.005 205.055 ;
        RECT 79.175 204.085 79.505 204.885 ;
        RECT 79.675 204.255 79.950 205.055 ;
        RECT 80.125 204.085 80.415 205.250 ;
        RECT 80.585 204.975 82.345 205.275 ;
        RECT 80.750 204.425 81.165 204.805 ;
        RECT 81.335 204.595 81.505 204.975 ;
        RECT 81.675 204.425 82.005 204.785 ;
        RECT 82.175 204.595 82.345 204.975 ;
        RECT 82.515 205.055 84.550 205.265 ;
        RECT 82.515 204.425 82.845 205.055 ;
        RECT 80.750 204.255 82.845 204.425 ;
        RECT 83.015 204.085 83.265 204.885 ;
        RECT 83.435 204.255 83.605 205.055 ;
        RECT 83.775 204.085 84.105 204.885 ;
        RECT 84.275 204.255 84.550 205.055 ;
        RECT 84.730 205.055 86.765 205.265 ;
        RECT 84.730 204.255 85.005 205.055 ;
        RECT 85.175 204.085 85.505 204.885 ;
        RECT 85.675 204.255 85.845 205.055 ;
        RECT 86.015 204.085 86.265 204.885 ;
        RECT 86.435 204.425 86.765 205.055 ;
        RECT 86.935 204.975 88.695 205.275 ;
        RECT 89.500 205.185 89.670 205.395 ;
        RECT 88.955 205.015 89.670 205.185 ;
        RECT 89.925 205.160 90.095 205.890 ;
        RECT 90.270 205.795 90.530 206.635 ;
        RECT 90.705 205.865 94.215 206.635 ;
        RECT 94.385 205.885 95.595 206.635 ;
        RECT 95.765 206.135 96.065 206.465 ;
        RECT 96.235 206.155 96.510 206.635 ;
        RECT 90.705 205.345 92.355 205.865 ;
        RECT 86.935 204.595 87.105 204.975 ;
        RECT 87.275 204.425 87.605 204.785 ;
        RECT 87.775 204.595 87.945 204.975 ;
        RECT 88.115 204.425 88.530 204.805 ;
        RECT 86.435 204.255 88.530 204.425 ;
        RECT 88.955 204.255 89.125 205.015 ;
        RECT 89.340 204.085 89.670 204.845 ;
        RECT 89.840 204.255 90.095 205.160 ;
        RECT 90.270 204.085 90.530 205.235 ;
        RECT 92.525 205.175 94.215 205.695 ;
        RECT 94.385 205.345 94.905 205.885 ;
        RECT 95.075 205.175 95.595 205.715 ;
        RECT 90.705 204.085 94.215 205.175 ;
        RECT 94.385 204.085 95.595 205.175 ;
        RECT 95.765 205.225 95.935 206.135 ;
        RECT 96.690 205.985 96.985 206.375 ;
        RECT 97.155 206.155 97.410 206.635 ;
        RECT 97.585 205.985 97.845 206.375 ;
        RECT 98.015 206.155 98.295 206.635 ;
        RECT 96.105 205.395 96.455 205.965 ;
        RECT 96.690 205.815 98.340 205.985 ;
        RECT 96.625 205.475 97.765 205.645 ;
        RECT 96.625 205.225 96.795 205.475 ;
        RECT 97.935 205.305 98.340 205.815 ;
        RECT 98.525 205.865 101.115 206.635 ;
        RECT 101.375 206.085 101.545 206.465 ;
        RECT 101.760 206.255 102.090 206.635 ;
        RECT 101.375 205.915 102.090 206.085 ;
        RECT 98.525 205.345 99.735 205.865 ;
        RECT 95.765 205.055 96.795 205.225 ;
        RECT 97.585 205.135 98.340 205.305 ;
        RECT 99.905 205.175 101.115 205.695 ;
        RECT 101.285 205.365 101.640 205.735 ;
        RECT 101.920 205.725 102.090 205.915 ;
        RECT 102.260 205.890 102.515 206.465 ;
        RECT 101.920 205.395 102.175 205.725 ;
        RECT 101.345 205.355 101.515 205.365 ;
        RECT 101.920 205.185 102.090 205.395 ;
        RECT 95.765 204.255 96.075 205.055 ;
        RECT 97.585 204.885 97.845 205.135 ;
        RECT 96.245 204.085 96.555 204.885 ;
        RECT 96.725 204.715 97.845 204.885 ;
        RECT 96.725 204.255 96.985 204.715 ;
        RECT 97.155 204.085 97.410 204.545 ;
        RECT 97.585 204.255 97.845 204.715 ;
        RECT 98.015 204.085 98.300 204.955 ;
        RECT 98.525 204.085 101.115 205.175 ;
        RECT 101.375 205.015 102.090 205.185 ;
        RECT 102.345 205.160 102.515 205.890 ;
        RECT 102.690 205.795 102.950 206.635 ;
        RECT 103.125 206.135 103.425 206.465 ;
        RECT 103.595 206.155 103.870 206.635 ;
        RECT 101.375 204.255 101.545 205.015 ;
        RECT 101.760 204.085 102.090 204.845 ;
        RECT 102.260 204.255 102.515 205.160 ;
        RECT 102.690 204.085 102.950 205.235 ;
        RECT 103.125 205.225 103.295 206.135 ;
        RECT 104.050 205.985 104.345 206.375 ;
        RECT 104.515 206.155 104.770 206.635 ;
        RECT 104.945 205.985 105.205 206.375 ;
        RECT 105.375 206.155 105.655 206.635 ;
        RECT 103.465 205.395 103.815 205.965 ;
        RECT 104.050 205.815 105.700 205.985 ;
        RECT 105.885 205.910 106.175 206.635 ;
        RECT 107.325 206.155 107.605 206.635 ;
        RECT 107.775 205.985 108.035 206.375 ;
        RECT 108.210 206.155 108.465 206.635 ;
        RECT 108.635 205.985 108.930 206.375 ;
        RECT 109.110 206.155 109.385 206.635 ;
        RECT 109.555 206.135 109.855 206.465 ;
        RECT 103.985 205.475 105.125 205.645 ;
        RECT 103.985 205.225 104.155 205.475 ;
        RECT 105.295 205.305 105.700 205.815 ;
        RECT 103.125 205.055 104.155 205.225 ;
        RECT 104.945 205.135 105.700 205.305 ;
        RECT 107.280 205.815 108.930 205.985 ;
        RECT 107.280 205.305 107.685 205.815 ;
        RECT 107.855 205.475 108.995 205.645 ;
        RECT 103.125 204.255 103.435 205.055 ;
        RECT 104.945 204.885 105.205 205.135 ;
        RECT 103.605 204.085 103.915 204.885 ;
        RECT 104.085 204.715 105.205 204.885 ;
        RECT 104.085 204.255 104.345 204.715 ;
        RECT 104.515 204.085 104.770 204.545 ;
        RECT 104.945 204.255 105.205 204.715 ;
        RECT 105.375 204.085 105.660 204.955 ;
        RECT 105.885 204.085 106.175 205.250 ;
        RECT 107.280 205.135 108.035 205.305 ;
        RECT 107.320 204.085 107.605 204.955 ;
        RECT 107.775 204.885 108.035 205.135 ;
        RECT 108.825 205.225 108.995 205.475 ;
        RECT 109.165 205.395 109.515 205.965 ;
        RECT 109.685 205.225 109.855 206.135 ;
        RECT 110.115 206.085 110.285 206.465 ;
        RECT 110.500 206.255 110.830 206.635 ;
        RECT 110.115 205.915 110.830 206.085 ;
        RECT 110.025 205.365 110.380 205.735 ;
        RECT 110.660 205.725 110.830 205.915 ;
        RECT 111.000 205.890 111.255 206.465 ;
        RECT 110.660 205.395 110.915 205.725 ;
        RECT 110.085 205.355 110.255 205.365 ;
        RECT 108.825 205.055 109.855 205.225 ;
        RECT 110.660 205.185 110.830 205.395 ;
        RECT 107.775 204.715 108.895 204.885 ;
        RECT 107.775 204.255 108.035 204.715 ;
        RECT 108.210 204.085 108.465 204.545 ;
        RECT 108.635 204.255 108.895 204.715 ;
        RECT 109.065 204.085 109.375 204.885 ;
        RECT 109.545 204.255 109.855 205.055 ;
        RECT 110.115 205.015 110.830 205.185 ;
        RECT 111.085 205.160 111.255 205.890 ;
        RECT 111.430 205.795 111.690 206.635 ;
        RECT 111.865 206.090 117.210 206.635 ;
        RECT 113.450 205.260 113.790 206.090 ;
        RECT 117.425 205.815 117.655 206.635 ;
        RECT 117.825 205.835 118.155 206.465 ;
        RECT 110.115 204.255 110.285 205.015 ;
        RECT 110.500 204.085 110.830 204.845 ;
        RECT 111.000 204.255 111.255 205.160 ;
        RECT 111.430 204.085 111.690 205.235 ;
        RECT 115.270 204.520 115.620 205.770 ;
        RECT 117.405 205.395 117.735 205.645 ;
        RECT 117.905 205.235 118.155 205.835 ;
        RECT 118.325 205.815 118.535 206.635 ;
        RECT 118.765 206.090 124.110 206.635 ;
        RECT 124.285 206.090 129.630 206.635 ;
        RECT 120.350 205.260 120.690 206.090 ;
        RECT 111.865 204.085 117.210 204.520 ;
        RECT 117.425 204.085 117.655 205.225 ;
        RECT 117.825 204.255 118.155 205.235 ;
        RECT 118.325 204.085 118.535 205.225 ;
        RECT 122.170 204.520 122.520 205.770 ;
        RECT 125.870 205.260 126.210 206.090 ;
        RECT 129.805 205.865 131.475 206.635 ;
        RECT 131.645 205.910 131.935 206.635 ;
        RECT 132.105 206.090 137.450 206.635 ;
        RECT 137.625 206.090 142.970 206.635 ;
        RECT 143.145 206.090 148.490 206.635 ;
        RECT 127.690 204.520 128.040 205.770 ;
        RECT 129.805 205.345 130.555 205.865 ;
        RECT 130.725 205.175 131.475 205.695 ;
        RECT 133.690 205.260 134.030 206.090 ;
        RECT 118.765 204.085 124.110 204.520 ;
        RECT 124.285 204.085 129.630 204.520 ;
        RECT 129.805 204.085 131.475 205.175 ;
        RECT 131.645 204.085 131.935 205.250 ;
        RECT 135.510 204.520 135.860 205.770 ;
        RECT 139.210 205.260 139.550 206.090 ;
        RECT 141.030 204.520 141.380 205.770 ;
        RECT 144.730 205.260 145.070 206.090 ;
        RECT 148.665 205.885 149.875 206.635 ;
        RECT 146.550 204.520 146.900 205.770 ;
        RECT 148.665 205.345 149.185 205.885 ;
        RECT 150.195 205.835 150.525 206.635 ;
        RECT 150.695 205.985 150.865 206.465 ;
        RECT 151.035 206.155 151.365 206.635 ;
        RECT 151.535 205.985 151.705 206.465 ;
        RECT 151.955 206.155 152.195 206.635 ;
        RECT 152.375 205.985 152.545 206.465 ;
        RECT 150.695 205.815 151.705 205.985 ;
        RECT 151.910 205.815 152.545 205.985 ;
        RECT 152.805 205.865 156.315 206.635 ;
        RECT 156.945 205.885 158.155 206.635 ;
        RECT 149.355 205.175 149.875 205.715 ;
        RECT 150.695 205.695 151.195 205.815 ;
        RECT 150.695 205.275 151.190 205.695 ;
        RECT 151.910 205.645 152.080 205.815 ;
        RECT 151.580 205.475 152.080 205.645 ;
        RECT 132.105 204.085 137.450 204.520 ;
        RECT 137.625 204.085 142.970 204.520 ;
        RECT 143.145 204.085 148.490 204.520 ;
        RECT 148.665 204.085 149.875 205.175 ;
        RECT 150.195 204.085 150.525 205.235 ;
        RECT 150.695 205.105 151.705 205.275 ;
        RECT 150.695 204.255 150.865 205.105 ;
        RECT 151.035 204.085 151.365 204.885 ;
        RECT 151.535 204.255 151.705 205.105 ;
        RECT 151.910 205.235 152.080 205.475 ;
        RECT 152.250 205.405 152.630 205.645 ;
        RECT 152.805 205.345 154.455 205.865 ;
        RECT 151.910 205.065 152.625 205.235 ;
        RECT 154.625 205.175 156.315 205.695 ;
        RECT 151.885 204.085 152.125 204.885 ;
        RECT 152.295 204.255 152.625 205.065 ;
        RECT 152.805 204.085 156.315 205.175 ;
        RECT 156.945 205.175 157.465 205.715 ;
        RECT 157.635 205.345 158.155 205.885 ;
        RECT 156.945 204.085 158.155 205.175 ;
        RECT 2.760 203.915 158.240 204.085 ;
        RECT 2.845 202.825 4.055 203.915 ;
        RECT 4.225 203.480 9.570 203.915 ;
        RECT 9.745 203.480 15.090 203.915 ;
        RECT 2.845 202.115 3.365 202.655 ;
        RECT 3.535 202.285 4.055 202.825 ;
        RECT 2.845 201.365 4.055 202.115 ;
        RECT 5.810 201.910 6.150 202.740 ;
        RECT 7.630 202.230 7.980 203.480 ;
        RECT 11.330 201.910 11.670 202.740 ;
        RECT 13.150 202.230 13.500 203.480 ;
        RECT 15.725 202.750 16.015 203.915 ;
        RECT 16.185 203.480 21.530 203.915 ;
        RECT 21.705 203.480 27.050 203.915 ;
        RECT 4.225 201.365 9.570 201.910 ;
        RECT 9.745 201.365 15.090 201.910 ;
        RECT 15.725 201.365 16.015 202.090 ;
        RECT 17.770 201.910 18.110 202.740 ;
        RECT 19.590 202.230 19.940 203.480 ;
        RECT 23.290 201.910 23.630 202.740 ;
        RECT 25.110 202.230 25.460 203.480 ;
        RECT 27.225 202.825 28.435 203.915 ;
        RECT 27.225 202.115 27.745 202.655 ;
        RECT 27.915 202.285 28.435 202.825 ;
        RECT 28.605 202.750 28.895 203.915 ;
        RECT 29.065 203.480 34.410 203.915 ;
        RECT 34.585 203.480 39.930 203.915 ;
        RECT 16.185 201.365 21.530 201.910 ;
        RECT 21.705 201.365 27.050 201.910 ;
        RECT 27.225 201.365 28.435 202.115 ;
        RECT 28.605 201.365 28.895 202.090 ;
        RECT 30.650 201.910 30.990 202.740 ;
        RECT 32.470 202.230 32.820 203.480 ;
        RECT 36.170 201.910 36.510 202.740 ;
        RECT 37.990 202.230 38.340 203.480 ;
        RECT 40.105 202.825 41.315 203.915 ;
        RECT 40.105 202.115 40.625 202.655 ;
        RECT 40.795 202.285 41.315 202.825 ;
        RECT 41.485 202.750 41.775 203.915 ;
        RECT 41.945 203.480 47.290 203.915 ;
        RECT 47.465 203.480 52.810 203.915 ;
        RECT 29.065 201.365 34.410 201.910 ;
        RECT 34.585 201.365 39.930 201.910 ;
        RECT 40.105 201.365 41.315 202.115 ;
        RECT 41.485 201.365 41.775 202.090 ;
        RECT 43.530 201.910 43.870 202.740 ;
        RECT 45.350 202.230 45.700 203.480 ;
        RECT 49.050 201.910 49.390 202.740 ;
        RECT 50.870 202.230 51.220 203.480 ;
        RECT 52.985 202.825 54.195 203.915 ;
        RECT 52.985 202.115 53.505 202.655 ;
        RECT 53.675 202.285 54.195 202.825 ;
        RECT 54.365 202.750 54.655 203.915 ;
        RECT 54.825 203.480 60.170 203.915 ;
        RECT 41.945 201.365 47.290 201.910 ;
        RECT 47.465 201.365 52.810 201.910 ;
        RECT 52.985 201.365 54.195 202.115 ;
        RECT 54.365 201.365 54.655 202.090 ;
        RECT 56.410 201.910 56.750 202.740 ;
        RECT 58.230 202.230 58.580 203.480 ;
        RECT 60.345 202.825 62.935 203.915 ;
        RECT 60.345 202.135 61.555 202.655 ;
        RECT 61.725 202.305 62.935 202.825 ;
        RECT 63.565 203.195 64.025 203.745 ;
        RECT 64.215 203.195 64.545 203.915 ;
        RECT 54.825 201.365 60.170 201.910 ;
        RECT 60.345 201.365 62.935 202.135 ;
        RECT 63.565 201.825 63.815 203.195 ;
        RECT 64.745 203.025 65.045 203.575 ;
        RECT 65.215 203.245 65.495 203.915 ;
        RECT 64.105 202.855 65.045 203.025 ;
        RECT 64.105 202.605 64.275 202.855 ;
        RECT 65.415 202.605 65.680 202.965 ;
        RECT 65.865 202.825 67.075 203.915 ;
        RECT 63.985 202.275 64.275 202.605 ;
        RECT 64.445 202.355 64.785 202.605 ;
        RECT 65.005 202.355 65.680 202.605 ;
        RECT 64.105 202.185 64.275 202.275 ;
        RECT 64.105 201.995 65.495 202.185 ;
        RECT 63.565 201.535 64.125 201.825 ;
        RECT 64.295 201.365 64.545 201.825 ;
        RECT 65.165 201.635 65.495 201.995 ;
        RECT 65.865 202.115 66.385 202.655 ;
        RECT 66.555 202.285 67.075 202.825 ;
        RECT 67.245 202.750 67.535 203.915 ;
        RECT 67.705 203.480 73.050 203.915 ;
        RECT 65.865 201.365 67.075 202.115 ;
        RECT 67.245 201.365 67.535 202.090 ;
        RECT 69.290 201.910 69.630 202.740 ;
        RECT 71.110 202.230 71.460 203.480 ;
        RECT 73.225 202.825 74.895 203.915 ;
        RECT 75.230 203.575 77.325 203.745 ;
        RECT 75.230 203.195 75.645 203.575 ;
        RECT 75.815 203.025 75.985 203.405 ;
        RECT 76.155 203.215 76.485 203.575 ;
        RECT 76.655 203.025 76.825 203.405 ;
        RECT 73.225 202.135 73.975 202.655 ;
        RECT 74.145 202.305 74.895 202.825 ;
        RECT 75.065 202.725 76.825 203.025 ;
        RECT 76.995 202.945 77.325 203.575 ;
        RECT 77.495 203.115 77.745 203.915 ;
        RECT 77.915 202.945 78.085 203.745 ;
        RECT 78.255 203.115 78.585 203.915 ;
        RECT 78.755 202.945 79.030 203.745 ;
        RECT 76.995 202.735 79.030 202.945 ;
        RECT 80.125 202.750 80.415 203.915 ;
        RECT 80.675 202.985 80.845 203.745 ;
        RECT 81.060 203.155 81.390 203.915 ;
        RECT 80.675 202.815 81.390 202.985 ;
        RECT 81.560 202.840 81.815 203.745 ;
        RECT 75.065 202.185 75.465 202.725 ;
        RECT 75.635 202.355 77.000 202.555 ;
        RECT 77.320 202.355 78.980 202.555 ;
        RECT 80.585 202.265 80.940 202.635 ;
        RECT 81.220 202.605 81.390 202.815 ;
        RECT 81.220 202.275 81.475 202.605 ;
        RECT 67.705 201.365 73.050 201.910 ;
        RECT 73.225 201.365 74.895 202.135 ;
        RECT 75.065 202.005 78.585 202.185 ;
        RECT 75.280 201.365 75.565 201.835 ;
        RECT 75.735 201.535 76.065 202.005 ;
        RECT 76.235 201.365 76.405 201.835 ;
        RECT 76.575 201.535 76.905 202.005 ;
        RECT 77.075 201.365 77.245 201.835 ;
        RECT 77.415 201.535 77.745 202.005 ;
        RECT 77.915 201.365 78.085 201.835 ;
        RECT 78.255 201.535 78.585 202.005 ;
        RECT 78.755 201.365 79.030 202.185 ;
        RECT 80.125 201.365 80.415 202.090 ;
        RECT 81.220 202.085 81.390 202.275 ;
        RECT 81.645 202.125 81.815 202.840 ;
        RECT 81.990 202.765 82.250 203.915 ;
        RECT 82.425 203.480 87.770 203.915 ;
        RECT 81.565 202.110 81.815 202.125 ;
        RECT 80.675 201.915 81.390 202.085 ;
        RECT 80.675 201.535 80.845 201.915 ;
        RECT 81.060 201.365 81.390 201.745 ;
        RECT 81.560 201.535 81.815 202.110 ;
        RECT 81.990 201.365 82.250 202.205 ;
        RECT 84.010 201.910 84.350 202.740 ;
        RECT 85.830 202.230 86.180 203.480 ;
        RECT 87.945 202.825 91.455 203.915 ;
        RECT 91.625 202.825 92.835 203.915 ;
        RECT 87.945 202.135 89.595 202.655 ;
        RECT 89.765 202.305 91.455 202.825 ;
        RECT 82.425 201.365 87.770 201.910 ;
        RECT 87.945 201.365 91.455 202.135 ;
        RECT 91.625 202.115 92.145 202.655 ;
        RECT 92.315 202.285 92.835 202.825 ;
        RECT 93.005 202.750 93.295 203.915 ;
        RECT 93.465 203.480 98.810 203.915 ;
        RECT 98.985 203.480 104.330 203.915 ;
        RECT 91.625 201.365 92.835 202.115 ;
        RECT 93.005 201.365 93.295 202.090 ;
        RECT 95.050 201.910 95.390 202.740 ;
        RECT 96.870 202.230 97.220 203.480 ;
        RECT 100.570 201.910 100.910 202.740 ;
        RECT 102.390 202.230 102.740 203.480 ;
        RECT 104.505 202.825 105.715 203.915 ;
        RECT 104.505 202.115 105.025 202.655 ;
        RECT 105.195 202.285 105.715 202.825 ;
        RECT 105.885 202.750 106.175 203.915 ;
        RECT 106.345 203.480 111.690 203.915 ;
        RECT 111.865 203.480 117.210 203.915 ;
        RECT 93.465 201.365 98.810 201.910 ;
        RECT 98.985 201.365 104.330 201.910 ;
        RECT 104.505 201.365 105.715 202.115 ;
        RECT 105.885 201.365 106.175 202.090 ;
        RECT 107.930 201.910 108.270 202.740 ;
        RECT 109.750 202.230 110.100 203.480 ;
        RECT 113.450 201.910 113.790 202.740 ;
        RECT 115.270 202.230 115.620 203.480 ;
        RECT 117.385 202.825 118.595 203.915 ;
        RECT 117.385 202.115 117.905 202.655 ;
        RECT 118.075 202.285 118.595 202.825 ;
        RECT 118.765 202.750 119.055 203.915 ;
        RECT 119.225 203.480 124.570 203.915 ;
        RECT 124.745 203.480 130.090 203.915 ;
        RECT 106.345 201.365 111.690 201.910 ;
        RECT 111.865 201.365 117.210 201.910 ;
        RECT 117.385 201.365 118.595 202.115 ;
        RECT 118.765 201.365 119.055 202.090 ;
        RECT 120.810 201.910 121.150 202.740 ;
        RECT 122.630 202.230 122.980 203.480 ;
        RECT 126.330 201.910 126.670 202.740 ;
        RECT 128.150 202.230 128.500 203.480 ;
        RECT 130.265 202.825 131.475 203.915 ;
        RECT 130.265 202.115 130.785 202.655 ;
        RECT 130.955 202.285 131.475 202.825 ;
        RECT 131.645 202.750 131.935 203.915 ;
        RECT 132.105 203.480 137.450 203.915 ;
        RECT 137.625 203.480 142.970 203.915 ;
        RECT 119.225 201.365 124.570 201.910 ;
        RECT 124.745 201.365 130.090 201.910 ;
        RECT 130.265 201.365 131.475 202.115 ;
        RECT 131.645 201.365 131.935 202.090 ;
        RECT 133.690 201.910 134.030 202.740 ;
        RECT 135.510 202.230 135.860 203.480 ;
        RECT 139.210 201.910 139.550 202.740 ;
        RECT 141.030 202.230 141.380 203.480 ;
        RECT 143.145 202.825 144.355 203.915 ;
        RECT 143.145 202.115 143.665 202.655 ;
        RECT 143.835 202.285 144.355 202.825 ;
        RECT 144.525 202.750 144.815 203.915 ;
        RECT 144.985 203.480 150.330 203.915 ;
        RECT 150.505 203.480 155.850 203.915 ;
        RECT 132.105 201.365 137.450 201.910 ;
        RECT 137.625 201.365 142.970 201.910 ;
        RECT 143.145 201.365 144.355 202.115 ;
        RECT 144.525 201.365 144.815 202.090 ;
        RECT 146.570 201.910 146.910 202.740 ;
        RECT 148.390 202.230 148.740 203.480 ;
        RECT 152.090 201.910 152.430 202.740 ;
        RECT 153.910 202.230 154.260 203.480 ;
        RECT 156.945 202.825 158.155 203.915 ;
        RECT 156.945 202.285 157.465 202.825 ;
        RECT 157.635 202.115 158.155 202.655 ;
        RECT 144.985 201.365 150.330 201.910 ;
        RECT 150.505 201.365 155.850 201.910 ;
        RECT 156.945 201.365 158.155 202.115 ;
        RECT 2.760 201.195 158.240 201.365 ;
        RECT 1.000 199.470 159.040 200.470 ;
        RECT 1.000 198.160 3.150 199.470 ;
        RECT 3.630 198.640 5.790 198.990 ;
        RECT 45.630 198.640 47.790 198.990 ;
        RECT 48.270 198.160 48.450 199.470 ;
        RECT 48.930 198.640 51.090 198.990 ;
        RECT 90.930 198.640 93.090 198.990 ;
        RECT 93.570 198.160 159.040 199.470 ;
        RECT 1.000 197.150 159.040 198.160 ;
        RECT 8.035 166.150 19.850 166.500 ;
        RECT 8.035 158.660 10.950 166.150 ;
        RECT 11.580 165.640 11.930 165.810 ;
        RECT 12.220 165.640 12.570 165.810 ;
        RECT 12.860 165.640 13.210 165.810 ;
        RECT 13.500 165.640 13.850 165.810 ;
        RECT 14.140 165.640 14.490 165.810 ;
        RECT 14.780 165.640 15.130 165.810 ;
        RECT 15.420 165.640 15.770 165.810 ;
        RECT 16.060 165.640 16.410 165.810 ;
        RECT 16.700 165.640 17.050 165.810 ;
        RECT 17.340 165.640 17.690 165.810 ;
        RECT 17.980 165.640 18.330 165.810 ;
        RECT 11.350 159.385 11.520 165.425 ;
        RECT 11.990 159.385 12.160 165.425 ;
        RECT 12.630 159.385 12.800 165.425 ;
        RECT 13.270 159.385 13.440 165.425 ;
        RECT 13.910 159.385 14.080 165.425 ;
        RECT 14.550 159.385 14.720 165.425 ;
        RECT 15.190 159.385 15.360 165.425 ;
        RECT 15.830 159.385 16.000 165.425 ;
        RECT 16.470 159.385 16.640 165.425 ;
        RECT 17.110 159.385 17.280 165.425 ;
        RECT 17.750 159.385 17.920 165.425 ;
        RECT 18.390 159.385 18.560 165.425 ;
        RECT 11.580 159.000 11.930 159.170 ;
        RECT 12.220 159.000 12.570 159.170 ;
        RECT 12.860 159.000 13.210 159.170 ;
        RECT 13.500 159.000 13.850 159.170 ;
        RECT 14.140 159.000 14.490 159.170 ;
        RECT 14.780 159.000 15.130 159.170 ;
        RECT 15.420 159.000 15.770 159.170 ;
        RECT 16.060 159.000 16.410 159.170 ;
        RECT 16.700 159.000 17.050 159.170 ;
        RECT 17.340 159.000 17.690 159.170 ;
        RECT 17.980 159.000 18.330 159.170 ;
        RECT 11.600 158.660 17.550 158.665 ;
        RECT 18.960 158.660 19.850 166.150 ;
        RECT 8.035 158.490 19.850 158.660 ;
        RECT 8.035 156.500 17.550 158.490 ;
        RECT 17.950 157.080 18.120 158.120 ;
        RECT 18.390 157.080 18.560 158.120 ;
        RECT 18.090 156.695 18.420 156.865 ;
        RECT 18.960 156.500 19.850 158.490 ;
        RECT 8.035 156.000 19.850 156.500 ;
        RECT 8.035 148.660 10.950 156.000 ;
        RECT 11.580 155.640 11.930 155.810 ;
        RECT 12.220 155.640 12.570 155.810 ;
        RECT 12.860 155.640 13.210 155.810 ;
        RECT 13.500 155.640 13.850 155.810 ;
        RECT 14.140 155.640 14.490 155.810 ;
        RECT 14.780 155.640 15.130 155.810 ;
        RECT 15.420 155.640 15.770 155.810 ;
        RECT 16.060 155.640 16.410 155.810 ;
        RECT 16.700 155.640 17.050 155.810 ;
        RECT 17.340 155.640 17.690 155.810 ;
        RECT 17.980 155.640 18.330 155.810 ;
        RECT 11.350 149.385 11.520 155.425 ;
        RECT 11.990 149.385 12.160 155.425 ;
        RECT 12.630 149.385 12.800 155.425 ;
        RECT 13.270 149.385 13.440 155.425 ;
        RECT 13.910 149.385 14.080 155.425 ;
        RECT 14.550 149.385 14.720 155.425 ;
        RECT 15.190 149.385 15.360 155.425 ;
        RECT 15.830 149.385 16.000 155.425 ;
        RECT 16.470 149.385 16.640 155.425 ;
        RECT 17.110 149.385 17.280 155.425 ;
        RECT 17.750 149.385 17.920 155.425 ;
        RECT 18.390 149.385 18.560 155.425 ;
        RECT 11.580 149.000 11.930 149.170 ;
        RECT 12.220 149.000 12.570 149.170 ;
        RECT 12.860 149.000 13.210 149.170 ;
        RECT 13.500 149.000 13.850 149.170 ;
        RECT 14.140 149.000 14.490 149.170 ;
        RECT 14.780 149.000 15.130 149.170 ;
        RECT 15.420 149.000 15.770 149.170 ;
        RECT 16.060 149.000 16.410 149.170 ;
        RECT 16.700 149.000 17.050 149.170 ;
        RECT 17.340 149.000 17.690 149.170 ;
        RECT 17.980 149.000 18.330 149.170 ;
        RECT 11.600 148.660 17.550 148.665 ;
        RECT 18.960 148.660 19.850 156.000 ;
        RECT 8.035 148.490 19.850 148.660 ;
        RECT 8.035 146.500 17.550 148.490 ;
        RECT 17.950 147.080 18.120 148.120 ;
        RECT 18.390 147.080 18.560 148.120 ;
        RECT 18.090 146.695 18.420 146.865 ;
        RECT 18.960 146.500 19.850 148.490 ;
        RECT 8.035 146.000 19.850 146.500 ;
        RECT 8.035 138.660 10.950 146.000 ;
        RECT 11.580 145.640 11.930 145.810 ;
        RECT 12.220 145.640 12.570 145.810 ;
        RECT 12.860 145.640 13.210 145.810 ;
        RECT 13.500 145.640 13.850 145.810 ;
        RECT 14.140 145.640 14.490 145.810 ;
        RECT 14.780 145.640 15.130 145.810 ;
        RECT 15.420 145.640 15.770 145.810 ;
        RECT 16.060 145.640 16.410 145.810 ;
        RECT 16.700 145.640 17.050 145.810 ;
        RECT 17.340 145.640 17.690 145.810 ;
        RECT 17.980 145.640 18.330 145.810 ;
        RECT 11.350 139.385 11.520 145.425 ;
        RECT 11.990 139.385 12.160 145.425 ;
        RECT 12.630 139.385 12.800 145.425 ;
        RECT 13.270 139.385 13.440 145.425 ;
        RECT 13.910 139.385 14.080 145.425 ;
        RECT 14.550 139.385 14.720 145.425 ;
        RECT 15.190 139.385 15.360 145.425 ;
        RECT 15.830 139.385 16.000 145.425 ;
        RECT 16.470 139.385 16.640 145.425 ;
        RECT 17.110 139.385 17.280 145.425 ;
        RECT 17.750 139.385 17.920 145.425 ;
        RECT 18.390 139.385 18.560 145.425 ;
        RECT 11.580 139.000 11.930 139.170 ;
        RECT 12.220 139.000 12.570 139.170 ;
        RECT 12.860 139.000 13.210 139.170 ;
        RECT 13.500 139.000 13.850 139.170 ;
        RECT 14.140 139.000 14.490 139.170 ;
        RECT 14.780 139.000 15.130 139.170 ;
        RECT 15.420 139.000 15.770 139.170 ;
        RECT 16.060 139.000 16.410 139.170 ;
        RECT 16.700 139.000 17.050 139.170 ;
        RECT 17.340 139.000 17.690 139.170 ;
        RECT 17.980 139.000 18.330 139.170 ;
        RECT 11.600 138.660 17.550 138.665 ;
        RECT 18.960 138.660 19.850 146.000 ;
        RECT 8.035 138.490 19.850 138.660 ;
        RECT 8.035 136.500 17.550 138.490 ;
        RECT 17.950 137.080 18.120 138.120 ;
        RECT 18.390 137.080 18.560 138.120 ;
        RECT 18.090 136.695 18.420 136.865 ;
        RECT 18.960 136.500 19.850 138.490 ;
        RECT 8.035 136.000 19.850 136.500 ;
        RECT 8.035 128.660 10.950 136.000 ;
        RECT 11.580 135.640 11.930 135.810 ;
        RECT 12.220 135.640 12.570 135.810 ;
        RECT 12.860 135.640 13.210 135.810 ;
        RECT 13.500 135.640 13.850 135.810 ;
        RECT 14.140 135.640 14.490 135.810 ;
        RECT 14.780 135.640 15.130 135.810 ;
        RECT 15.420 135.640 15.770 135.810 ;
        RECT 16.060 135.640 16.410 135.810 ;
        RECT 16.700 135.640 17.050 135.810 ;
        RECT 17.340 135.640 17.690 135.810 ;
        RECT 17.980 135.640 18.330 135.810 ;
        RECT 11.350 129.385 11.520 135.425 ;
        RECT 11.990 129.385 12.160 135.425 ;
        RECT 12.630 129.385 12.800 135.425 ;
        RECT 13.270 129.385 13.440 135.425 ;
        RECT 13.910 129.385 14.080 135.425 ;
        RECT 14.550 129.385 14.720 135.425 ;
        RECT 15.190 129.385 15.360 135.425 ;
        RECT 15.830 129.385 16.000 135.425 ;
        RECT 16.470 129.385 16.640 135.425 ;
        RECT 17.110 129.385 17.280 135.425 ;
        RECT 17.750 129.385 17.920 135.425 ;
        RECT 18.390 129.385 18.560 135.425 ;
        RECT 11.580 129.000 11.930 129.170 ;
        RECT 12.220 129.000 12.570 129.170 ;
        RECT 12.860 129.000 13.210 129.170 ;
        RECT 13.500 129.000 13.850 129.170 ;
        RECT 14.140 129.000 14.490 129.170 ;
        RECT 14.780 129.000 15.130 129.170 ;
        RECT 15.420 129.000 15.770 129.170 ;
        RECT 16.060 129.000 16.410 129.170 ;
        RECT 16.700 129.000 17.050 129.170 ;
        RECT 17.340 129.000 17.690 129.170 ;
        RECT 17.980 129.000 18.330 129.170 ;
        RECT 11.600 128.660 17.550 128.665 ;
        RECT 18.960 128.660 19.850 136.000 ;
        RECT 8.035 128.490 19.850 128.660 ;
        RECT 8.035 126.500 17.550 128.490 ;
        RECT 17.950 127.080 18.120 128.120 ;
        RECT 18.390 127.080 18.560 128.120 ;
        RECT 18.090 126.695 18.420 126.865 ;
        RECT 18.960 126.500 19.850 128.490 ;
        RECT 8.035 126.000 19.850 126.500 ;
        RECT 8.035 118.660 10.950 126.000 ;
        RECT 11.580 125.640 11.930 125.810 ;
        RECT 12.220 125.640 12.570 125.810 ;
        RECT 12.860 125.640 13.210 125.810 ;
        RECT 13.500 125.640 13.850 125.810 ;
        RECT 14.140 125.640 14.490 125.810 ;
        RECT 14.780 125.640 15.130 125.810 ;
        RECT 15.420 125.640 15.770 125.810 ;
        RECT 16.060 125.640 16.410 125.810 ;
        RECT 16.700 125.640 17.050 125.810 ;
        RECT 17.340 125.640 17.690 125.810 ;
        RECT 17.980 125.640 18.330 125.810 ;
        RECT 11.350 119.385 11.520 125.425 ;
        RECT 11.990 119.385 12.160 125.425 ;
        RECT 12.630 119.385 12.800 125.425 ;
        RECT 13.270 119.385 13.440 125.425 ;
        RECT 13.910 119.385 14.080 125.425 ;
        RECT 14.550 119.385 14.720 125.425 ;
        RECT 15.190 119.385 15.360 125.425 ;
        RECT 15.830 119.385 16.000 125.425 ;
        RECT 16.470 119.385 16.640 125.425 ;
        RECT 17.110 119.385 17.280 125.425 ;
        RECT 17.750 119.385 17.920 125.425 ;
        RECT 18.390 119.385 18.560 125.425 ;
        RECT 11.580 119.000 11.930 119.170 ;
        RECT 12.220 119.000 12.570 119.170 ;
        RECT 12.860 119.000 13.210 119.170 ;
        RECT 13.500 119.000 13.850 119.170 ;
        RECT 14.140 119.000 14.490 119.170 ;
        RECT 14.780 119.000 15.130 119.170 ;
        RECT 15.420 119.000 15.770 119.170 ;
        RECT 16.060 119.000 16.410 119.170 ;
        RECT 16.700 119.000 17.050 119.170 ;
        RECT 17.340 119.000 17.690 119.170 ;
        RECT 17.980 119.000 18.330 119.170 ;
        RECT 11.600 118.660 17.550 118.665 ;
        RECT 18.960 118.660 19.850 126.000 ;
        RECT 8.035 118.490 19.850 118.660 ;
        RECT 8.035 116.500 17.550 118.490 ;
        RECT 17.950 117.080 18.120 118.120 ;
        RECT 18.390 117.080 18.560 118.120 ;
        RECT 18.090 116.695 18.420 116.865 ;
        RECT 18.960 116.500 19.850 118.490 ;
        RECT 8.035 116.000 19.850 116.500 ;
        RECT 8.035 108.660 10.950 116.000 ;
        RECT 11.580 115.640 11.930 115.810 ;
        RECT 12.220 115.640 12.570 115.810 ;
        RECT 12.860 115.640 13.210 115.810 ;
        RECT 13.500 115.640 13.850 115.810 ;
        RECT 14.140 115.640 14.490 115.810 ;
        RECT 14.780 115.640 15.130 115.810 ;
        RECT 15.420 115.640 15.770 115.810 ;
        RECT 16.060 115.640 16.410 115.810 ;
        RECT 16.700 115.640 17.050 115.810 ;
        RECT 17.340 115.640 17.690 115.810 ;
        RECT 17.980 115.640 18.330 115.810 ;
        RECT 11.350 109.385 11.520 115.425 ;
        RECT 11.990 109.385 12.160 115.425 ;
        RECT 12.630 109.385 12.800 115.425 ;
        RECT 13.270 109.385 13.440 115.425 ;
        RECT 13.910 109.385 14.080 115.425 ;
        RECT 14.550 109.385 14.720 115.425 ;
        RECT 15.190 109.385 15.360 115.425 ;
        RECT 15.830 109.385 16.000 115.425 ;
        RECT 16.470 109.385 16.640 115.425 ;
        RECT 17.110 109.385 17.280 115.425 ;
        RECT 17.750 109.385 17.920 115.425 ;
        RECT 18.390 109.385 18.560 115.425 ;
        RECT 11.580 109.000 11.930 109.170 ;
        RECT 12.220 109.000 12.570 109.170 ;
        RECT 12.860 109.000 13.210 109.170 ;
        RECT 13.500 109.000 13.850 109.170 ;
        RECT 14.140 109.000 14.490 109.170 ;
        RECT 14.780 109.000 15.130 109.170 ;
        RECT 15.420 109.000 15.770 109.170 ;
        RECT 16.060 109.000 16.410 109.170 ;
        RECT 16.700 109.000 17.050 109.170 ;
        RECT 17.340 109.000 17.690 109.170 ;
        RECT 17.980 109.000 18.330 109.170 ;
        RECT 11.600 108.660 17.550 108.665 ;
        RECT 18.960 108.660 19.850 116.000 ;
        RECT 8.035 108.490 19.850 108.660 ;
        RECT 8.035 106.500 17.550 108.490 ;
        RECT 17.950 107.080 18.120 108.120 ;
        RECT 18.390 107.080 18.560 108.120 ;
        RECT 18.090 106.695 18.420 106.865 ;
        RECT 18.960 106.500 19.850 108.490 ;
        RECT 8.035 106.000 19.850 106.500 ;
        RECT 8.035 98.660 10.950 106.000 ;
        RECT 11.580 105.640 11.930 105.810 ;
        RECT 12.220 105.640 12.570 105.810 ;
        RECT 12.860 105.640 13.210 105.810 ;
        RECT 13.500 105.640 13.850 105.810 ;
        RECT 14.140 105.640 14.490 105.810 ;
        RECT 14.780 105.640 15.130 105.810 ;
        RECT 15.420 105.640 15.770 105.810 ;
        RECT 16.060 105.640 16.410 105.810 ;
        RECT 16.700 105.640 17.050 105.810 ;
        RECT 17.340 105.640 17.690 105.810 ;
        RECT 17.980 105.640 18.330 105.810 ;
        RECT 11.350 99.385 11.520 105.425 ;
        RECT 11.990 99.385 12.160 105.425 ;
        RECT 12.630 99.385 12.800 105.425 ;
        RECT 13.270 99.385 13.440 105.425 ;
        RECT 13.910 99.385 14.080 105.425 ;
        RECT 14.550 99.385 14.720 105.425 ;
        RECT 15.190 99.385 15.360 105.425 ;
        RECT 15.830 99.385 16.000 105.425 ;
        RECT 16.470 99.385 16.640 105.425 ;
        RECT 17.110 99.385 17.280 105.425 ;
        RECT 17.750 99.385 17.920 105.425 ;
        RECT 18.390 99.385 18.560 105.425 ;
        RECT 11.580 99.000 11.930 99.170 ;
        RECT 12.220 99.000 12.570 99.170 ;
        RECT 12.860 99.000 13.210 99.170 ;
        RECT 13.500 99.000 13.850 99.170 ;
        RECT 14.140 99.000 14.490 99.170 ;
        RECT 14.780 99.000 15.130 99.170 ;
        RECT 15.420 99.000 15.770 99.170 ;
        RECT 16.060 99.000 16.410 99.170 ;
        RECT 16.700 99.000 17.050 99.170 ;
        RECT 17.340 99.000 17.690 99.170 ;
        RECT 17.980 99.000 18.330 99.170 ;
        RECT 11.600 98.660 17.550 98.665 ;
        RECT 18.960 98.660 19.850 106.000 ;
        RECT 8.035 98.490 19.850 98.660 ;
        RECT 8.035 96.500 17.550 98.490 ;
        RECT 17.950 97.080 18.120 98.120 ;
        RECT 18.390 97.080 18.560 98.120 ;
        RECT 18.090 96.695 18.420 96.865 ;
        RECT 18.960 96.500 19.850 98.490 ;
        RECT 8.035 96.000 19.850 96.500 ;
        RECT 8.035 88.660 10.950 96.000 ;
        RECT 11.580 95.640 11.930 95.810 ;
        RECT 12.220 95.640 12.570 95.810 ;
        RECT 12.860 95.640 13.210 95.810 ;
        RECT 13.500 95.640 13.850 95.810 ;
        RECT 14.140 95.640 14.490 95.810 ;
        RECT 14.780 95.640 15.130 95.810 ;
        RECT 15.420 95.640 15.770 95.810 ;
        RECT 16.060 95.640 16.410 95.810 ;
        RECT 16.700 95.640 17.050 95.810 ;
        RECT 17.340 95.640 17.690 95.810 ;
        RECT 17.980 95.640 18.330 95.810 ;
        RECT 11.350 89.385 11.520 95.425 ;
        RECT 11.990 89.385 12.160 95.425 ;
        RECT 12.630 89.385 12.800 95.425 ;
        RECT 13.270 89.385 13.440 95.425 ;
        RECT 13.910 89.385 14.080 95.425 ;
        RECT 14.550 89.385 14.720 95.425 ;
        RECT 15.190 89.385 15.360 95.425 ;
        RECT 15.830 89.385 16.000 95.425 ;
        RECT 16.470 89.385 16.640 95.425 ;
        RECT 17.110 89.385 17.280 95.425 ;
        RECT 17.750 89.385 17.920 95.425 ;
        RECT 18.390 89.385 18.560 95.425 ;
        RECT 11.580 89.000 11.930 89.170 ;
        RECT 12.220 89.000 12.570 89.170 ;
        RECT 12.860 89.000 13.210 89.170 ;
        RECT 13.500 89.000 13.850 89.170 ;
        RECT 14.140 89.000 14.490 89.170 ;
        RECT 14.780 89.000 15.130 89.170 ;
        RECT 15.420 89.000 15.770 89.170 ;
        RECT 16.060 89.000 16.410 89.170 ;
        RECT 16.700 89.000 17.050 89.170 ;
        RECT 17.340 89.000 17.690 89.170 ;
        RECT 17.980 89.000 18.330 89.170 ;
        RECT 11.600 88.660 17.550 88.665 ;
        RECT 18.960 88.660 19.850 96.000 ;
        RECT 8.035 88.490 19.850 88.660 ;
        RECT 8.035 86.500 17.550 88.490 ;
        RECT 17.950 87.080 18.120 88.120 ;
        RECT 18.390 87.080 18.560 88.120 ;
        RECT 18.090 86.695 18.420 86.865 ;
        RECT 18.960 86.500 19.850 88.490 ;
        RECT 8.035 86.000 19.850 86.500 ;
        RECT 8.035 78.660 10.950 86.000 ;
        RECT 11.580 85.640 11.930 85.810 ;
        RECT 12.220 85.640 12.570 85.810 ;
        RECT 12.860 85.640 13.210 85.810 ;
        RECT 13.500 85.640 13.850 85.810 ;
        RECT 14.140 85.640 14.490 85.810 ;
        RECT 14.780 85.640 15.130 85.810 ;
        RECT 15.420 85.640 15.770 85.810 ;
        RECT 16.060 85.640 16.410 85.810 ;
        RECT 16.700 85.640 17.050 85.810 ;
        RECT 17.340 85.640 17.690 85.810 ;
        RECT 17.980 85.640 18.330 85.810 ;
        RECT 11.350 79.385 11.520 85.425 ;
        RECT 11.990 79.385 12.160 85.425 ;
        RECT 12.630 79.385 12.800 85.425 ;
        RECT 13.270 79.385 13.440 85.425 ;
        RECT 13.910 79.385 14.080 85.425 ;
        RECT 14.550 79.385 14.720 85.425 ;
        RECT 15.190 79.385 15.360 85.425 ;
        RECT 15.830 79.385 16.000 85.425 ;
        RECT 16.470 79.385 16.640 85.425 ;
        RECT 17.110 79.385 17.280 85.425 ;
        RECT 17.750 79.385 17.920 85.425 ;
        RECT 18.390 79.385 18.560 85.425 ;
        RECT 11.580 79.000 11.930 79.170 ;
        RECT 12.220 79.000 12.570 79.170 ;
        RECT 12.860 79.000 13.210 79.170 ;
        RECT 13.500 79.000 13.850 79.170 ;
        RECT 14.140 79.000 14.490 79.170 ;
        RECT 14.780 79.000 15.130 79.170 ;
        RECT 15.420 79.000 15.770 79.170 ;
        RECT 16.060 79.000 16.410 79.170 ;
        RECT 16.700 79.000 17.050 79.170 ;
        RECT 17.340 79.000 17.690 79.170 ;
        RECT 17.980 79.000 18.330 79.170 ;
        RECT 11.600 78.660 17.550 78.665 ;
        RECT 18.960 78.660 19.850 86.000 ;
        RECT 8.035 78.490 19.850 78.660 ;
        RECT 8.035 76.500 17.550 78.490 ;
        RECT 17.950 77.080 18.120 78.120 ;
        RECT 18.390 77.080 18.560 78.120 ;
        RECT 18.090 76.695 18.420 76.865 ;
        RECT 18.960 76.500 19.850 78.490 ;
        RECT 8.035 76.000 19.850 76.500 ;
        RECT 8.035 68.660 10.950 76.000 ;
        RECT 11.580 75.640 11.930 75.810 ;
        RECT 12.220 75.640 12.570 75.810 ;
        RECT 12.860 75.640 13.210 75.810 ;
        RECT 13.500 75.640 13.850 75.810 ;
        RECT 14.140 75.640 14.490 75.810 ;
        RECT 14.780 75.640 15.130 75.810 ;
        RECT 15.420 75.640 15.770 75.810 ;
        RECT 16.060 75.640 16.410 75.810 ;
        RECT 16.700 75.640 17.050 75.810 ;
        RECT 17.340 75.640 17.690 75.810 ;
        RECT 17.980 75.640 18.330 75.810 ;
        RECT 11.350 69.385 11.520 75.425 ;
        RECT 11.990 69.385 12.160 75.425 ;
        RECT 12.630 69.385 12.800 75.425 ;
        RECT 13.270 69.385 13.440 75.425 ;
        RECT 13.910 69.385 14.080 75.425 ;
        RECT 14.550 69.385 14.720 75.425 ;
        RECT 15.190 69.385 15.360 75.425 ;
        RECT 15.830 69.385 16.000 75.425 ;
        RECT 16.470 69.385 16.640 75.425 ;
        RECT 17.110 69.385 17.280 75.425 ;
        RECT 17.750 69.385 17.920 75.425 ;
        RECT 18.390 69.385 18.560 75.425 ;
        RECT 11.580 69.000 11.930 69.170 ;
        RECT 12.220 69.000 12.570 69.170 ;
        RECT 12.860 69.000 13.210 69.170 ;
        RECT 13.500 69.000 13.850 69.170 ;
        RECT 14.140 69.000 14.490 69.170 ;
        RECT 14.780 69.000 15.130 69.170 ;
        RECT 15.420 69.000 15.770 69.170 ;
        RECT 16.060 69.000 16.410 69.170 ;
        RECT 16.700 69.000 17.050 69.170 ;
        RECT 17.340 69.000 17.690 69.170 ;
        RECT 17.980 69.000 18.330 69.170 ;
        RECT 11.600 68.660 17.550 68.665 ;
        RECT 18.960 68.660 19.850 76.000 ;
        RECT 8.035 68.490 19.850 68.660 ;
        RECT 8.035 66.500 17.550 68.490 ;
        RECT 17.950 67.080 18.120 68.120 ;
        RECT 18.390 67.080 18.560 68.120 ;
        RECT 18.090 66.695 18.420 66.865 ;
        RECT 18.960 66.500 19.850 68.490 ;
        RECT 8.035 66.000 19.850 66.500 ;
        RECT 8.035 58.660 10.950 66.000 ;
        RECT 11.580 65.640 11.930 65.810 ;
        RECT 12.220 65.640 12.570 65.810 ;
        RECT 12.860 65.640 13.210 65.810 ;
        RECT 13.500 65.640 13.850 65.810 ;
        RECT 14.140 65.640 14.490 65.810 ;
        RECT 14.780 65.640 15.130 65.810 ;
        RECT 15.420 65.640 15.770 65.810 ;
        RECT 16.060 65.640 16.410 65.810 ;
        RECT 16.700 65.640 17.050 65.810 ;
        RECT 17.340 65.640 17.690 65.810 ;
        RECT 17.980 65.640 18.330 65.810 ;
        RECT 11.350 59.385 11.520 65.425 ;
        RECT 11.990 59.385 12.160 65.425 ;
        RECT 12.630 59.385 12.800 65.425 ;
        RECT 13.270 59.385 13.440 65.425 ;
        RECT 13.910 59.385 14.080 65.425 ;
        RECT 14.550 59.385 14.720 65.425 ;
        RECT 15.190 59.385 15.360 65.425 ;
        RECT 15.830 59.385 16.000 65.425 ;
        RECT 16.470 59.385 16.640 65.425 ;
        RECT 17.110 59.385 17.280 65.425 ;
        RECT 17.750 59.385 17.920 65.425 ;
        RECT 18.390 59.385 18.560 65.425 ;
        RECT 11.580 59.000 11.930 59.170 ;
        RECT 12.220 59.000 12.570 59.170 ;
        RECT 12.860 59.000 13.210 59.170 ;
        RECT 13.500 59.000 13.850 59.170 ;
        RECT 14.140 59.000 14.490 59.170 ;
        RECT 14.780 59.000 15.130 59.170 ;
        RECT 15.420 59.000 15.770 59.170 ;
        RECT 16.060 59.000 16.410 59.170 ;
        RECT 16.700 59.000 17.050 59.170 ;
        RECT 17.340 59.000 17.690 59.170 ;
        RECT 17.980 59.000 18.330 59.170 ;
        RECT 11.600 58.660 17.550 58.665 ;
        RECT 18.960 58.660 19.850 66.000 ;
        RECT 8.035 58.490 19.850 58.660 ;
        RECT 8.035 56.500 17.550 58.490 ;
        RECT 17.950 57.080 18.120 58.120 ;
        RECT 18.390 57.080 18.560 58.120 ;
        RECT 18.090 56.695 18.420 56.865 ;
        RECT 18.960 56.500 19.850 58.490 ;
        RECT 8.035 56.000 19.850 56.500 ;
        RECT 8.035 48.660 10.950 56.000 ;
        RECT 11.580 55.640 11.930 55.810 ;
        RECT 12.220 55.640 12.570 55.810 ;
        RECT 12.860 55.640 13.210 55.810 ;
        RECT 13.500 55.640 13.850 55.810 ;
        RECT 14.140 55.640 14.490 55.810 ;
        RECT 14.780 55.640 15.130 55.810 ;
        RECT 15.420 55.640 15.770 55.810 ;
        RECT 16.060 55.640 16.410 55.810 ;
        RECT 16.700 55.640 17.050 55.810 ;
        RECT 17.340 55.640 17.690 55.810 ;
        RECT 17.980 55.640 18.330 55.810 ;
        RECT 11.350 49.385 11.520 55.425 ;
        RECT 11.990 49.385 12.160 55.425 ;
        RECT 12.630 49.385 12.800 55.425 ;
        RECT 13.270 49.385 13.440 55.425 ;
        RECT 13.910 49.385 14.080 55.425 ;
        RECT 14.550 49.385 14.720 55.425 ;
        RECT 15.190 49.385 15.360 55.425 ;
        RECT 15.830 49.385 16.000 55.425 ;
        RECT 16.470 49.385 16.640 55.425 ;
        RECT 17.110 49.385 17.280 55.425 ;
        RECT 17.750 49.385 17.920 55.425 ;
        RECT 18.390 49.385 18.560 55.425 ;
        RECT 11.580 49.000 11.930 49.170 ;
        RECT 12.220 49.000 12.570 49.170 ;
        RECT 12.860 49.000 13.210 49.170 ;
        RECT 13.500 49.000 13.850 49.170 ;
        RECT 14.140 49.000 14.490 49.170 ;
        RECT 14.780 49.000 15.130 49.170 ;
        RECT 15.420 49.000 15.770 49.170 ;
        RECT 16.060 49.000 16.410 49.170 ;
        RECT 16.700 49.000 17.050 49.170 ;
        RECT 17.340 49.000 17.690 49.170 ;
        RECT 17.980 49.000 18.330 49.170 ;
        RECT 11.600 48.660 17.550 48.665 ;
        RECT 18.960 48.660 19.850 56.000 ;
        RECT 8.035 48.490 19.850 48.660 ;
        RECT 8.035 46.500 17.550 48.490 ;
        RECT 17.950 47.080 18.120 48.120 ;
        RECT 18.390 47.080 18.560 48.120 ;
        RECT 18.090 46.695 18.420 46.865 ;
        RECT 18.960 46.500 19.850 48.490 ;
        RECT 8.035 46.000 19.850 46.500 ;
        RECT 8.035 38.660 10.950 46.000 ;
        RECT 11.580 45.640 11.930 45.810 ;
        RECT 12.220 45.640 12.570 45.810 ;
        RECT 12.860 45.640 13.210 45.810 ;
        RECT 13.500 45.640 13.850 45.810 ;
        RECT 14.140 45.640 14.490 45.810 ;
        RECT 14.780 45.640 15.130 45.810 ;
        RECT 15.420 45.640 15.770 45.810 ;
        RECT 16.060 45.640 16.410 45.810 ;
        RECT 16.700 45.640 17.050 45.810 ;
        RECT 17.340 45.640 17.690 45.810 ;
        RECT 17.980 45.640 18.330 45.810 ;
        RECT 11.350 39.385 11.520 45.425 ;
        RECT 11.990 39.385 12.160 45.425 ;
        RECT 12.630 39.385 12.800 45.425 ;
        RECT 13.270 39.385 13.440 45.425 ;
        RECT 13.910 39.385 14.080 45.425 ;
        RECT 14.550 39.385 14.720 45.425 ;
        RECT 15.190 39.385 15.360 45.425 ;
        RECT 15.830 39.385 16.000 45.425 ;
        RECT 16.470 39.385 16.640 45.425 ;
        RECT 17.110 39.385 17.280 45.425 ;
        RECT 17.750 39.385 17.920 45.425 ;
        RECT 18.390 39.385 18.560 45.425 ;
        RECT 11.580 39.000 11.930 39.170 ;
        RECT 12.220 39.000 12.570 39.170 ;
        RECT 12.860 39.000 13.210 39.170 ;
        RECT 13.500 39.000 13.850 39.170 ;
        RECT 14.140 39.000 14.490 39.170 ;
        RECT 14.780 39.000 15.130 39.170 ;
        RECT 15.420 39.000 15.770 39.170 ;
        RECT 16.060 39.000 16.410 39.170 ;
        RECT 16.700 39.000 17.050 39.170 ;
        RECT 17.340 39.000 17.690 39.170 ;
        RECT 17.980 39.000 18.330 39.170 ;
        RECT 11.600 38.660 17.550 38.665 ;
        RECT 18.960 38.660 19.850 46.000 ;
        RECT 8.035 38.490 19.850 38.660 ;
        RECT 8.035 36.500 17.550 38.490 ;
        RECT 17.950 37.080 18.120 38.120 ;
        RECT 18.390 37.080 18.560 38.120 ;
        RECT 18.090 36.695 18.420 36.865 ;
        RECT 18.960 36.500 19.850 38.490 ;
        RECT 8.035 36.000 19.850 36.500 ;
        RECT 8.035 28.660 10.950 36.000 ;
        RECT 11.580 35.640 11.930 35.810 ;
        RECT 12.220 35.640 12.570 35.810 ;
        RECT 12.860 35.640 13.210 35.810 ;
        RECT 13.500 35.640 13.850 35.810 ;
        RECT 14.140 35.640 14.490 35.810 ;
        RECT 14.780 35.640 15.130 35.810 ;
        RECT 15.420 35.640 15.770 35.810 ;
        RECT 16.060 35.640 16.410 35.810 ;
        RECT 16.700 35.640 17.050 35.810 ;
        RECT 17.340 35.640 17.690 35.810 ;
        RECT 17.980 35.640 18.330 35.810 ;
        RECT 11.350 29.385 11.520 35.425 ;
        RECT 11.990 29.385 12.160 35.425 ;
        RECT 12.630 29.385 12.800 35.425 ;
        RECT 13.270 29.385 13.440 35.425 ;
        RECT 13.910 29.385 14.080 35.425 ;
        RECT 14.550 29.385 14.720 35.425 ;
        RECT 15.190 29.385 15.360 35.425 ;
        RECT 15.830 29.385 16.000 35.425 ;
        RECT 16.470 29.385 16.640 35.425 ;
        RECT 17.110 29.385 17.280 35.425 ;
        RECT 17.750 29.385 17.920 35.425 ;
        RECT 18.390 29.385 18.560 35.425 ;
        RECT 11.580 29.000 11.930 29.170 ;
        RECT 12.220 29.000 12.570 29.170 ;
        RECT 12.860 29.000 13.210 29.170 ;
        RECT 13.500 29.000 13.850 29.170 ;
        RECT 14.140 29.000 14.490 29.170 ;
        RECT 14.780 29.000 15.130 29.170 ;
        RECT 15.420 29.000 15.770 29.170 ;
        RECT 16.060 29.000 16.410 29.170 ;
        RECT 16.700 29.000 17.050 29.170 ;
        RECT 17.340 29.000 17.690 29.170 ;
        RECT 17.980 29.000 18.330 29.170 ;
        RECT 11.600 28.660 17.550 28.665 ;
        RECT 18.960 28.660 19.850 36.000 ;
        RECT 8.035 28.490 19.850 28.660 ;
        RECT 8.035 26.500 17.550 28.490 ;
        RECT 17.950 27.080 18.120 28.120 ;
        RECT 18.390 27.080 18.560 28.120 ;
        RECT 18.090 26.695 18.420 26.865 ;
        RECT 18.960 26.500 19.850 28.490 ;
        RECT 8.035 26.000 19.850 26.500 ;
        RECT 8.035 18.660 10.950 26.000 ;
        RECT 11.580 25.640 11.930 25.810 ;
        RECT 12.220 25.640 12.570 25.810 ;
        RECT 12.860 25.640 13.210 25.810 ;
        RECT 13.500 25.640 13.850 25.810 ;
        RECT 14.140 25.640 14.490 25.810 ;
        RECT 14.780 25.640 15.130 25.810 ;
        RECT 15.420 25.640 15.770 25.810 ;
        RECT 16.060 25.640 16.410 25.810 ;
        RECT 16.700 25.640 17.050 25.810 ;
        RECT 17.340 25.640 17.690 25.810 ;
        RECT 17.980 25.640 18.330 25.810 ;
        RECT 11.350 19.385 11.520 25.425 ;
        RECT 11.990 19.385 12.160 25.425 ;
        RECT 12.630 19.385 12.800 25.425 ;
        RECT 13.270 19.385 13.440 25.425 ;
        RECT 13.910 19.385 14.080 25.425 ;
        RECT 14.550 19.385 14.720 25.425 ;
        RECT 15.190 19.385 15.360 25.425 ;
        RECT 15.830 19.385 16.000 25.425 ;
        RECT 16.470 19.385 16.640 25.425 ;
        RECT 17.110 19.385 17.280 25.425 ;
        RECT 17.750 19.385 17.920 25.425 ;
        RECT 18.390 19.385 18.560 25.425 ;
        RECT 11.580 19.000 11.930 19.170 ;
        RECT 12.220 19.000 12.570 19.170 ;
        RECT 12.860 19.000 13.210 19.170 ;
        RECT 13.500 19.000 13.850 19.170 ;
        RECT 14.140 19.000 14.490 19.170 ;
        RECT 14.780 19.000 15.130 19.170 ;
        RECT 15.420 19.000 15.770 19.170 ;
        RECT 16.060 19.000 16.410 19.170 ;
        RECT 16.700 19.000 17.050 19.170 ;
        RECT 17.340 19.000 17.690 19.170 ;
        RECT 17.980 19.000 18.330 19.170 ;
        RECT 11.600 18.660 17.550 18.665 ;
        RECT 18.960 18.660 19.850 26.000 ;
        RECT 8.035 18.490 19.850 18.660 ;
        RECT 8.035 16.500 17.550 18.490 ;
        RECT 17.950 17.080 18.120 18.120 ;
        RECT 18.390 17.080 18.560 18.120 ;
        RECT 18.090 16.695 18.420 16.865 ;
        RECT 18.960 16.500 19.850 18.490 ;
        RECT 8.035 16.000 19.850 16.500 ;
        RECT 8.035 8.660 10.950 16.000 ;
        RECT 11.580 15.640 11.930 15.810 ;
        RECT 12.220 15.640 12.570 15.810 ;
        RECT 12.860 15.640 13.210 15.810 ;
        RECT 13.500 15.640 13.850 15.810 ;
        RECT 14.140 15.640 14.490 15.810 ;
        RECT 14.780 15.640 15.130 15.810 ;
        RECT 15.420 15.640 15.770 15.810 ;
        RECT 16.060 15.640 16.410 15.810 ;
        RECT 16.700 15.640 17.050 15.810 ;
        RECT 17.340 15.640 17.690 15.810 ;
        RECT 17.980 15.640 18.330 15.810 ;
        RECT 11.350 9.385 11.520 15.425 ;
        RECT 11.990 9.385 12.160 15.425 ;
        RECT 12.630 9.385 12.800 15.425 ;
        RECT 13.270 9.385 13.440 15.425 ;
        RECT 13.910 9.385 14.080 15.425 ;
        RECT 14.550 9.385 14.720 15.425 ;
        RECT 15.190 9.385 15.360 15.425 ;
        RECT 15.830 9.385 16.000 15.425 ;
        RECT 16.470 9.385 16.640 15.425 ;
        RECT 17.110 9.385 17.280 15.425 ;
        RECT 17.750 9.385 17.920 15.425 ;
        RECT 18.390 9.385 18.560 15.425 ;
        RECT 11.580 9.000 11.930 9.170 ;
        RECT 12.220 9.000 12.570 9.170 ;
        RECT 12.860 9.000 13.210 9.170 ;
        RECT 13.500 9.000 13.850 9.170 ;
        RECT 14.140 9.000 14.490 9.170 ;
        RECT 14.780 9.000 15.130 9.170 ;
        RECT 15.420 9.000 15.770 9.170 ;
        RECT 16.060 9.000 16.410 9.170 ;
        RECT 16.700 9.000 17.050 9.170 ;
        RECT 17.340 9.000 17.690 9.170 ;
        RECT 17.980 9.000 18.330 9.170 ;
        RECT 11.600 8.660 17.550 8.665 ;
        RECT 18.960 8.660 19.850 16.000 ;
        RECT 8.035 8.490 19.850 8.660 ;
        RECT 8.035 6.350 17.550 8.490 ;
        RECT 17.950 7.080 18.120 8.120 ;
        RECT 18.390 7.080 18.560 8.120 ;
        RECT 18.090 6.695 18.420 6.865 ;
        RECT 18.960 6.350 19.850 8.490 ;
        RECT 8.035 6.000 19.850 6.350 ;
        RECT 20.025 164.060 26.350 166.500 ;
        RECT 20.025 158.660 20.910 164.060 ;
        RECT 21.540 163.550 21.890 163.720 ;
        RECT 22.180 163.550 22.530 163.720 ;
        RECT 22.820 163.550 23.170 163.720 ;
        RECT 23.460 163.550 23.810 163.720 ;
        RECT 24.100 163.550 24.450 163.720 ;
        RECT 21.310 159.340 21.480 163.380 ;
        RECT 21.950 159.340 22.120 163.380 ;
        RECT 22.590 159.340 22.760 163.380 ;
        RECT 23.230 159.340 23.400 163.380 ;
        RECT 23.870 159.340 24.040 163.380 ;
        RECT 24.510 159.340 24.680 163.380 ;
        RECT 21.540 159.000 21.890 159.170 ;
        RECT 22.180 159.000 22.530 159.170 ;
        RECT 22.820 159.000 23.170 159.170 ;
        RECT 23.460 159.000 23.810 159.170 ;
        RECT 24.100 159.000 24.450 159.170 ;
        RECT 22.325 158.660 23.450 158.665 ;
        RECT 25.080 158.660 26.350 164.060 ;
        RECT 20.025 158.460 26.350 158.660 ;
        RECT 20.025 156.500 20.910 158.460 ;
        RECT 22.320 158.450 26.350 158.460 ;
        RECT 21.310 157.050 21.480 158.090 ;
        RECT 21.750 157.050 21.920 158.090 ;
        RECT 21.450 156.710 21.780 156.880 ;
        RECT 22.320 156.500 23.550 158.450 ;
        RECT 23.950 157.040 24.120 158.080 ;
        RECT 24.390 157.040 24.560 158.080 ;
        RECT 24.090 156.700 24.420 156.870 ;
        RECT 24.960 156.500 26.350 158.450 ;
        RECT 20.025 154.060 26.350 156.500 ;
        RECT 20.025 148.660 20.910 154.060 ;
        RECT 21.540 153.550 21.890 153.720 ;
        RECT 22.180 153.550 22.530 153.720 ;
        RECT 22.820 153.550 23.170 153.720 ;
        RECT 23.460 153.550 23.810 153.720 ;
        RECT 24.100 153.550 24.450 153.720 ;
        RECT 21.310 149.340 21.480 153.380 ;
        RECT 21.950 149.340 22.120 153.380 ;
        RECT 22.590 149.340 22.760 153.380 ;
        RECT 23.230 149.340 23.400 153.380 ;
        RECT 23.870 149.340 24.040 153.380 ;
        RECT 24.510 149.340 24.680 153.380 ;
        RECT 21.540 149.000 21.890 149.170 ;
        RECT 22.180 149.000 22.530 149.170 ;
        RECT 22.820 149.000 23.170 149.170 ;
        RECT 23.460 149.000 23.810 149.170 ;
        RECT 24.100 149.000 24.450 149.170 ;
        RECT 22.325 148.660 23.450 148.665 ;
        RECT 25.080 148.660 26.350 154.060 ;
        RECT 20.025 148.460 26.350 148.660 ;
        RECT 20.025 146.500 20.910 148.460 ;
        RECT 22.320 148.450 26.350 148.460 ;
        RECT 21.310 147.050 21.480 148.090 ;
        RECT 21.750 147.050 21.920 148.090 ;
        RECT 21.450 146.710 21.780 146.880 ;
        RECT 22.320 146.500 23.550 148.450 ;
        RECT 23.950 147.040 24.120 148.080 ;
        RECT 24.390 147.040 24.560 148.080 ;
        RECT 24.090 146.700 24.420 146.870 ;
        RECT 24.960 146.500 26.350 148.450 ;
        RECT 20.025 144.060 26.350 146.500 ;
        RECT 20.025 138.660 20.910 144.060 ;
        RECT 21.540 143.550 21.890 143.720 ;
        RECT 22.180 143.550 22.530 143.720 ;
        RECT 22.820 143.550 23.170 143.720 ;
        RECT 23.460 143.550 23.810 143.720 ;
        RECT 24.100 143.550 24.450 143.720 ;
        RECT 21.310 139.340 21.480 143.380 ;
        RECT 21.950 139.340 22.120 143.380 ;
        RECT 22.590 139.340 22.760 143.380 ;
        RECT 23.230 139.340 23.400 143.380 ;
        RECT 23.870 139.340 24.040 143.380 ;
        RECT 24.510 139.340 24.680 143.380 ;
        RECT 21.540 139.000 21.890 139.170 ;
        RECT 22.180 139.000 22.530 139.170 ;
        RECT 22.820 139.000 23.170 139.170 ;
        RECT 23.460 139.000 23.810 139.170 ;
        RECT 24.100 139.000 24.450 139.170 ;
        RECT 22.325 138.660 23.450 138.665 ;
        RECT 25.080 138.660 26.350 144.060 ;
        RECT 20.025 138.460 26.350 138.660 ;
        RECT 20.025 136.500 20.910 138.460 ;
        RECT 22.320 138.450 26.350 138.460 ;
        RECT 21.310 137.050 21.480 138.090 ;
        RECT 21.750 137.050 21.920 138.090 ;
        RECT 21.450 136.710 21.780 136.880 ;
        RECT 22.320 136.500 23.550 138.450 ;
        RECT 23.950 137.040 24.120 138.080 ;
        RECT 24.390 137.040 24.560 138.080 ;
        RECT 24.090 136.700 24.420 136.870 ;
        RECT 24.960 136.500 26.350 138.450 ;
        RECT 20.025 134.060 26.350 136.500 ;
        RECT 20.025 128.660 20.910 134.060 ;
        RECT 21.540 133.550 21.890 133.720 ;
        RECT 22.180 133.550 22.530 133.720 ;
        RECT 22.820 133.550 23.170 133.720 ;
        RECT 23.460 133.550 23.810 133.720 ;
        RECT 24.100 133.550 24.450 133.720 ;
        RECT 21.310 129.340 21.480 133.380 ;
        RECT 21.950 129.340 22.120 133.380 ;
        RECT 22.590 129.340 22.760 133.380 ;
        RECT 23.230 129.340 23.400 133.380 ;
        RECT 23.870 129.340 24.040 133.380 ;
        RECT 24.510 129.340 24.680 133.380 ;
        RECT 21.540 129.000 21.890 129.170 ;
        RECT 22.180 129.000 22.530 129.170 ;
        RECT 22.820 129.000 23.170 129.170 ;
        RECT 23.460 129.000 23.810 129.170 ;
        RECT 24.100 129.000 24.450 129.170 ;
        RECT 22.325 128.660 23.450 128.665 ;
        RECT 25.080 128.660 26.350 134.060 ;
        RECT 20.025 128.460 26.350 128.660 ;
        RECT 20.025 126.500 20.910 128.460 ;
        RECT 22.320 128.450 26.350 128.460 ;
        RECT 21.310 127.050 21.480 128.090 ;
        RECT 21.750 127.050 21.920 128.090 ;
        RECT 21.450 126.710 21.780 126.880 ;
        RECT 22.320 126.500 23.550 128.450 ;
        RECT 23.950 127.040 24.120 128.080 ;
        RECT 24.390 127.040 24.560 128.080 ;
        RECT 24.090 126.700 24.420 126.870 ;
        RECT 24.960 126.500 26.350 128.450 ;
        RECT 20.025 124.060 26.350 126.500 ;
        RECT 20.025 118.660 20.910 124.060 ;
        RECT 21.540 123.550 21.890 123.720 ;
        RECT 22.180 123.550 22.530 123.720 ;
        RECT 22.820 123.550 23.170 123.720 ;
        RECT 23.460 123.550 23.810 123.720 ;
        RECT 24.100 123.550 24.450 123.720 ;
        RECT 21.310 119.340 21.480 123.380 ;
        RECT 21.950 119.340 22.120 123.380 ;
        RECT 22.590 119.340 22.760 123.380 ;
        RECT 23.230 119.340 23.400 123.380 ;
        RECT 23.870 119.340 24.040 123.380 ;
        RECT 24.510 119.340 24.680 123.380 ;
        RECT 21.540 119.000 21.890 119.170 ;
        RECT 22.180 119.000 22.530 119.170 ;
        RECT 22.820 119.000 23.170 119.170 ;
        RECT 23.460 119.000 23.810 119.170 ;
        RECT 24.100 119.000 24.450 119.170 ;
        RECT 22.325 118.660 23.450 118.665 ;
        RECT 25.080 118.660 26.350 124.060 ;
        RECT 20.025 118.460 26.350 118.660 ;
        RECT 20.025 116.500 20.910 118.460 ;
        RECT 22.320 118.450 26.350 118.460 ;
        RECT 21.310 117.050 21.480 118.090 ;
        RECT 21.750 117.050 21.920 118.090 ;
        RECT 21.450 116.710 21.780 116.880 ;
        RECT 22.320 116.500 23.550 118.450 ;
        RECT 23.950 117.040 24.120 118.080 ;
        RECT 24.390 117.040 24.560 118.080 ;
        RECT 24.090 116.700 24.420 116.870 ;
        RECT 24.960 116.500 26.350 118.450 ;
        RECT 20.025 114.060 26.350 116.500 ;
        RECT 20.025 108.660 20.910 114.060 ;
        RECT 21.540 113.550 21.890 113.720 ;
        RECT 22.180 113.550 22.530 113.720 ;
        RECT 22.820 113.550 23.170 113.720 ;
        RECT 23.460 113.550 23.810 113.720 ;
        RECT 24.100 113.550 24.450 113.720 ;
        RECT 21.310 109.340 21.480 113.380 ;
        RECT 21.950 109.340 22.120 113.380 ;
        RECT 22.590 109.340 22.760 113.380 ;
        RECT 23.230 109.340 23.400 113.380 ;
        RECT 23.870 109.340 24.040 113.380 ;
        RECT 24.510 109.340 24.680 113.380 ;
        RECT 21.540 109.000 21.890 109.170 ;
        RECT 22.180 109.000 22.530 109.170 ;
        RECT 22.820 109.000 23.170 109.170 ;
        RECT 23.460 109.000 23.810 109.170 ;
        RECT 24.100 109.000 24.450 109.170 ;
        RECT 22.325 108.660 23.450 108.665 ;
        RECT 25.080 108.660 26.350 114.060 ;
        RECT 20.025 108.460 26.350 108.660 ;
        RECT 20.025 106.500 20.910 108.460 ;
        RECT 22.320 108.450 26.350 108.460 ;
        RECT 21.310 107.050 21.480 108.090 ;
        RECT 21.750 107.050 21.920 108.090 ;
        RECT 21.450 106.710 21.780 106.880 ;
        RECT 22.320 106.500 23.550 108.450 ;
        RECT 23.950 107.040 24.120 108.080 ;
        RECT 24.390 107.040 24.560 108.080 ;
        RECT 24.090 106.700 24.420 106.870 ;
        RECT 24.960 106.500 26.350 108.450 ;
        RECT 20.025 104.060 26.350 106.500 ;
        RECT 20.025 98.660 20.910 104.060 ;
        RECT 21.540 103.550 21.890 103.720 ;
        RECT 22.180 103.550 22.530 103.720 ;
        RECT 22.820 103.550 23.170 103.720 ;
        RECT 23.460 103.550 23.810 103.720 ;
        RECT 24.100 103.550 24.450 103.720 ;
        RECT 21.310 99.340 21.480 103.380 ;
        RECT 21.950 99.340 22.120 103.380 ;
        RECT 22.590 99.340 22.760 103.380 ;
        RECT 23.230 99.340 23.400 103.380 ;
        RECT 23.870 99.340 24.040 103.380 ;
        RECT 24.510 99.340 24.680 103.380 ;
        RECT 21.540 99.000 21.890 99.170 ;
        RECT 22.180 99.000 22.530 99.170 ;
        RECT 22.820 99.000 23.170 99.170 ;
        RECT 23.460 99.000 23.810 99.170 ;
        RECT 24.100 99.000 24.450 99.170 ;
        RECT 22.325 98.660 23.450 98.665 ;
        RECT 25.080 98.660 26.350 104.060 ;
        RECT 20.025 98.460 26.350 98.660 ;
        RECT 20.025 96.500 20.910 98.460 ;
        RECT 22.320 98.450 26.350 98.460 ;
        RECT 21.310 97.050 21.480 98.090 ;
        RECT 21.750 97.050 21.920 98.090 ;
        RECT 21.450 96.710 21.780 96.880 ;
        RECT 22.320 96.500 23.550 98.450 ;
        RECT 23.950 97.040 24.120 98.080 ;
        RECT 24.390 97.040 24.560 98.080 ;
        RECT 24.090 96.700 24.420 96.870 ;
        RECT 24.960 96.500 26.350 98.450 ;
        RECT 20.025 94.060 26.350 96.500 ;
        RECT 20.025 88.660 20.910 94.060 ;
        RECT 21.540 93.550 21.890 93.720 ;
        RECT 22.180 93.550 22.530 93.720 ;
        RECT 22.820 93.550 23.170 93.720 ;
        RECT 23.460 93.550 23.810 93.720 ;
        RECT 24.100 93.550 24.450 93.720 ;
        RECT 21.310 89.340 21.480 93.380 ;
        RECT 21.950 89.340 22.120 93.380 ;
        RECT 22.590 89.340 22.760 93.380 ;
        RECT 23.230 89.340 23.400 93.380 ;
        RECT 23.870 89.340 24.040 93.380 ;
        RECT 24.510 89.340 24.680 93.380 ;
        RECT 21.540 89.000 21.890 89.170 ;
        RECT 22.180 89.000 22.530 89.170 ;
        RECT 22.820 89.000 23.170 89.170 ;
        RECT 23.460 89.000 23.810 89.170 ;
        RECT 24.100 89.000 24.450 89.170 ;
        RECT 22.325 88.660 23.450 88.665 ;
        RECT 25.080 88.660 26.350 94.060 ;
        RECT 20.025 88.460 26.350 88.660 ;
        RECT 20.025 86.500 20.910 88.460 ;
        RECT 22.320 88.450 26.350 88.460 ;
        RECT 21.310 87.050 21.480 88.090 ;
        RECT 21.750 87.050 21.920 88.090 ;
        RECT 21.450 86.710 21.780 86.880 ;
        RECT 22.320 86.500 23.550 88.450 ;
        RECT 23.950 87.040 24.120 88.080 ;
        RECT 24.390 87.040 24.560 88.080 ;
        RECT 24.090 86.700 24.420 86.870 ;
        RECT 24.960 86.500 26.350 88.450 ;
        RECT 20.025 84.060 26.350 86.500 ;
        RECT 20.025 78.660 20.910 84.060 ;
        RECT 21.540 83.550 21.890 83.720 ;
        RECT 22.180 83.550 22.530 83.720 ;
        RECT 22.820 83.550 23.170 83.720 ;
        RECT 23.460 83.550 23.810 83.720 ;
        RECT 24.100 83.550 24.450 83.720 ;
        RECT 21.310 79.340 21.480 83.380 ;
        RECT 21.950 79.340 22.120 83.380 ;
        RECT 22.590 79.340 22.760 83.380 ;
        RECT 23.230 79.340 23.400 83.380 ;
        RECT 23.870 79.340 24.040 83.380 ;
        RECT 24.510 79.340 24.680 83.380 ;
        RECT 21.540 79.000 21.890 79.170 ;
        RECT 22.180 79.000 22.530 79.170 ;
        RECT 22.820 79.000 23.170 79.170 ;
        RECT 23.460 79.000 23.810 79.170 ;
        RECT 24.100 79.000 24.450 79.170 ;
        RECT 22.325 78.660 23.450 78.665 ;
        RECT 25.080 78.660 26.350 84.060 ;
        RECT 20.025 78.460 26.350 78.660 ;
        RECT 20.025 76.500 20.910 78.460 ;
        RECT 22.320 78.450 26.350 78.460 ;
        RECT 21.310 77.050 21.480 78.090 ;
        RECT 21.750 77.050 21.920 78.090 ;
        RECT 21.450 76.710 21.780 76.880 ;
        RECT 22.320 76.500 23.550 78.450 ;
        RECT 23.950 77.040 24.120 78.080 ;
        RECT 24.390 77.040 24.560 78.080 ;
        RECT 24.090 76.700 24.420 76.870 ;
        RECT 24.960 76.500 26.350 78.450 ;
        RECT 20.025 74.060 26.350 76.500 ;
        RECT 20.025 68.660 20.910 74.060 ;
        RECT 21.540 73.550 21.890 73.720 ;
        RECT 22.180 73.550 22.530 73.720 ;
        RECT 22.820 73.550 23.170 73.720 ;
        RECT 23.460 73.550 23.810 73.720 ;
        RECT 24.100 73.550 24.450 73.720 ;
        RECT 21.310 69.340 21.480 73.380 ;
        RECT 21.950 69.340 22.120 73.380 ;
        RECT 22.590 69.340 22.760 73.380 ;
        RECT 23.230 69.340 23.400 73.380 ;
        RECT 23.870 69.340 24.040 73.380 ;
        RECT 24.510 69.340 24.680 73.380 ;
        RECT 21.540 69.000 21.890 69.170 ;
        RECT 22.180 69.000 22.530 69.170 ;
        RECT 22.820 69.000 23.170 69.170 ;
        RECT 23.460 69.000 23.810 69.170 ;
        RECT 24.100 69.000 24.450 69.170 ;
        RECT 22.325 68.660 23.450 68.665 ;
        RECT 25.080 68.660 26.350 74.060 ;
        RECT 20.025 68.460 26.350 68.660 ;
        RECT 20.025 66.500 20.910 68.460 ;
        RECT 22.320 68.450 26.350 68.460 ;
        RECT 21.310 67.050 21.480 68.090 ;
        RECT 21.750 67.050 21.920 68.090 ;
        RECT 21.450 66.710 21.780 66.880 ;
        RECT 22.320 66.500 23.550 68.450 ;
        RECT 23.950 67.040 24.120 68.080 ;
        RECT 24.390 67.040 24.560 68.080 ;
        RECT 24.090 66.700 24.420 66.870 ;
        RECT 24.960 66.500 26.350 68.450 ;
        RECT 20.025 64.060 26.350 66.500 ;
        RECT 20.025 58.660 20.910 64.060 ;
        RECT 21.540 63.550 21.890 63.720 ;
        RECT 22.180 63.550 22.530 63.720 ;
        RECT 22.820 63.550 23.170 63.720 ;
        RECT 23.460 63.550 23.810 63.720 ;
        RECT 24.100 63.550 24.450 63.720 ;
        RECT 21.310 59.340 21.480 63.380 ;
        RECT 21.950 59.340 22.120 63.380 ;
        RECT 22.590 59.340 22.760 63.380 ;
        RECT 23.230 59.340 23.400 63.380 ;
        RECT 23.870 59.340 24.040 63.380 ;
        RECT 24.510 59.340 24.680 63.380 ;
        RECT 21.540 59.000 21.890 59.170 ;
        RECT 22.180 59.000 22.530 59.170 ;
        RECT 22.820 59.000 23.170 59.170 ;
        RECT 23.460 59.000 23.810 59.170 ;
        RECT 24.100 59.000 24.450 59.170 ;
        RECT 22.325 58.660 23.450 58.665 ;
        RECT 25.080 58.660 26.350 64.060 ;
        RECT 20.025 58.460 26.350 58.660 ;
        RECT 20.025 56.500 20.910 58.460 ;
        RECT 22.320 58.450 26.350 58.460 ;
        RECT 21.310 57.050 21.480 58.090 ;
        RECT 21.750 57.050 21.920 58.090 ;
        RECT 21.450 56.710 21.780 56.880 ;
        RECT 22.320 56.500 23.550 58.450 ;
        RECT 23.950 57.040 24.120 58.080 ;
        RECT 24.390 57.040 24.560 58.080 ;
        RECT 24.090 56.700 24.420 56.870 ;
        RECT 24.960 56.500 26.350 58.450 ;
        RECT 20.025 54.060 26.350 56.500 ;
        RECT 20.025 48.660 20.910 54.060 ;
        RECT 21.540 53.550 21.890 53.720 ;
        RECT 22.180 53.550 22.530 53.720 ;
        RECT 22.820 53.550 23.170 53.720 ;
        RECT 23.460 53.550 23.810 53.720 ;
        RECT 24.100 53.550 24.450 53.720 ;
        RECT 21.310 49.340 21.480 53.380 ;
        RECT 21.950 49.340 22.120 53.380 ;
        RECT 22.590 49.340 22.760 53.380 ;
        RECT 23.230 49.340 23.400 53.380 ;
        RECT 23.870 49.340 24.040 53.380 ;
        RECT 24.510 49.340 24.680 53.380 ;
        RECT 21.540 49.000 21.890 49.170 ;
        RECT 22.180 49.000 22.530 49.170 ;
        RECT 22.820 49.000 23.170 49.170 ;
        RECT 23.460 49.000 23.810 49.170 ;
        RECT 24.100 49.000 24.450 49.170 ;
        RECT 22.325 48.660 23.450 48.665 ;
        RECT 25.080 48.660 26.350 54.060 ;
        RECT 20.025 48.460 26.350 48.660 ;
        RECT 20.025 46.500 20.910 48.460 ;
        RECT 22.320 48.450 26.350 48.460 ;
        RECT 21.310 47.050 21.480 48.090 ;
        RECT 21.750 47.050 21.920 48.090 ;
        RECT 21.450 46.710 21.780 46.880 ;
        RECT 22.320 46.500 23.550 48.450 ;
        RECT 23.950 47.040 24.120 48.080 ;
        RECT 24.390 47.040 24.560 48.080 ;
        RECT 24.090 46.700 24.420 46.870 ;
        RECT 24.960 46.500 26.350 48.450 ;
        RECT 20.025 44.060 26.350 46.500 ;
        RECT 20.025 38.660 20.910 44.060 ;
        RECT 21.540 43.550 21.890 43.720 ;
        RECT 22.180 43.550 22.530 43.720 ;
        RECT 22.820 43.550 23.170 43.720 ;
        RECT 23.460 43.550 23.810 43.720 ;
        RECT 24.100 43.550 24.450 43.720 ;
        RECT 21.310 39.340 21.480 43.380 ;
        RECT 21.950 39.340 22.120 43.380 ;
        RECT 22.590 39.340 22.760 43.380 ;
        RECT 23.230 39.340 23.400 43.380 ;
        RECT 23.870 39.340 24.040 43.380 ;
        RECT 24.510 39.340 24.680 43.380 ;
        RECT 21.540 39.000 21.890 39.170 ;
        RECT 22.180 39.000 22.530 39.170 ;
        RECT 22.820 39.000 23.170 39.170 ;
        RECT 23.460 39.000 23.810 39.170 ;
        RECT 24.100 39.000 24.450 39.170 ;
        RECT 22.325 38.660 23.450 38.665 ;
        RECT 25.080 38.660 26.350 44.060 ;
        RECT 20.025 38.460 26.350 38.660 ;
        RECT 20.025 36.500 20.910 38.460 ;
        RECT 22.320 38.450 26.350 38.460 ;
        RECT 21.310 37.050 21.480 38.090 ;
        RECT 21.750 37.050 21.920 38.090 ;
        RECT 21.450 36.710 21.780 36.880 ;
        RECT 22.320 36.500 23.550 38.450 ;
        RECT 23.950 37.040 24.120 38.080 ;
        RECT 24.390 37.040 24.560 38.080 ;
        RECT 24.090 36.700 24.420 36.870 ;
        RECT 24.960 36.500 26.350 38.450 ;
        RECT 20.025 34.060 26.350 36.500 ;
        RECT 20.025 28.660 20.910 34.060 ;
        RECT 21.540 33.550 21.890 33.720 ;
        RECT 22.180 33.550 22.530 33.720 ;
        RECT 22.820 33.550 23.170 33.720 ;
        RECT 23.460 33.550 23.810 33.720 ;
        RECT 24.100 33.550 24.450 33.720 ;
        RECT 21.310 29.340 21.480 33.380 ;
        RECT 21.950 29.340 22.120 33.380 ;
        RECT 22.590 29.340 22.760 33.380 ;
        RECT 23.230 29.340 23.400 33.380 ;
        RECT 23.870 29.340 24.040 33.380 ;
        RECT 24.510 29.340 24.680 33.380 ;
        RECT 21.540 29.000 21.890 29.170 ;
        RECT 22.180 29.000 22.530 29.170 ;
        RECT 22.820 29.000 23.170 29.170 ;
        RECT 23.460 29.000 23.810 29.170 ;
        RECT 24.100 29.000 24.450 29.170 ;
        RECT 22.325 28.660 23.450 28.665 ;
        RECT 25.080 28.660 26.350 34.060 ;
        RECT 20.025 28.460 26.350 28.660 ;
        RECT 20.025 26.500 20.910 28.460 ;
        RECT 22.320 28.450 26.350 28.460 ;
        RECT 21.310 27.050 21.480 28.090 ;
        RECT 21.750 27.050 21.920 28.090 ;
        RECT 21.450 26.710 21.780 26.880 ;
        RECT 22.320 26.500 23.550 28.450 ;
        RECT 23.950 27.040 24.120 28.080 ;
        RECT 24.390 27.040 24.560 28.080 ;
        RECT 24.090 26.700 24.420 26.870 ;
        RECT 24.960 26.500 26.350 28.450 ;
        RECT 20.025 24.060 26.350 26.500 ;
        RECT 20.025 18.660 20.910 24.060 ;
        RECT 21.540 23.550 21.890 23.720 ;
        RECT 22.180 23.550 22.530 23.720 ;
        RECT 22.820 23.550 23.170 23.720 ;
        RECT 23.460 23.550 23.810 23.720 ;
        RECT 24.100 23.550 24.450 23.720 ;
        RECT 21.310 19.340 21.480 23.380 ;
        RECT 21.950 19.340 22.120 23.380 ;
        RECT 22.590 19.340 22.760 23.380 ;
        RECT 23.230 19.340 23.400 23.380 ;
        RECT 23.870 19.340 24.040 23.380 ;
        RECT 24.510 19.340 24.680 23.380 ;
        RECT 21.540 19.000 21.890 19.170 ;
        RECT 22.180 19.000 22.530 19.170 ;
        RECT 22.820 19.000 23.170 19.170 ;
        RECT 23.460 19.000 23.810 19.170 ;
        RECT 24.100 19.000 24.450 19.170 ;
        RECT 22.325 18.660 23.450 18.665 ;
        RECT 25.080 18.660 26.350 24.060 ;
        RECT 20.025 18.460 26.350 18.660 ;
        RECT 20.025 16.500 20.910 18.460 ;
        RECT 22.320 18.450 26.350 18.460 ;
        RECT 21.310 17.050 21.480 18.090 ;
        RECT 21.750 17.050 21.920 18.090 ;
        RECT 21.450 16.710 21.780 16.880 ;
        RECT 22.320 16.500 23.550 18.450 ;
        RECT 23.950 17.040 24.120 18.080 ;
        RECT 24.390 17.040 24.560 18.080 ;
        RECT 24.090 16.700 24.420 16.870 ;
        RECT 24.960 16.500 26.350 18.450 ;
        RECT 20.025 14.060 26.350 16.500 ;
        RECT 20.025 8.660 20.910 14.060 ;
        RECT 21.540 13.550 21.890 13.720 ;
        RECT 22.180 13.550 22.530 13.720 ;
        RECT 22.820 13.550 23.170 13.720 ;
        RECT 23.460 13.550 23.810 13.720 ;
        RECT 24.100 13.550 24.450 13.720 ;
        RECT 21.310 9.340 21.480 13.380 ;
        RECT 21.950 9.340 22.120 13.380 ;
        RECT 22.590 9.340 22.760 13.380 ;
        RECT 23.230 9.340 23.400 13.380 ;
        RECT 23.870 9.340 24.040 13.380 ;
        RECT 24.510 9.340 24.680 13.380 ;
        RECT 21.540 9.000 21.890 9.170 ;
        RECT 22.180 9.000 22.530 9.170 ;
        RECT 22.820 9.000 23.170 9.170 ;
        RECT 23.460 9.000 23.810 9.170 ;
        RECT 24.100 9.000 24.450 9.170 ;
        RECT 22.325 8.660 23.450 8.665 ;
        RECT 25.080 8.660 26.350 14.060 ;
        RECT 20.025 8.460 26.350 8.660 ;
        RECT 20.025 6.370 20.910 8.460 ;
        RECT 22.320 8.450 26.350 8.460 ;
        RECT 21.310 7.050 21.480 8.090 ;
        RECT 21.750 7.050 21.920 8.090 ;
        RECT 21.450 6.710 21.780 6.880 ;
        RECT 22.320 6.370 23.550 8.450 ;
        RECT 23.950 7.040 24.120 8.080 ;
        RECT 24.390 7.040 24.560 8.080 ;
        RECT 24.090 6.700 24.420 6.870 ;
        RECT 20.025 6.360 23.550 6.370 ;
        RECT 24.960 6.360 26.350 8.450 ;
        RECT 20.025 6.000 26.350 6.360 ;
        RECT 133.640 166.140 143.390 166.490 ;
        RECT 133.640 158.650 134.490 166.140 ;
        RECT 135.120 165.630 135.470 165.800 ;
        RECT 135.760 165.630 136.110 165.800 ;
        RECT 136.400 165.630 136.750 165.800 ;
        RECT 137.040 165.630 137.390 165.800 ;
        RECT 137.680 165.630 138.030 165.800 ;
        RECT 138.320 165.630 138.670 165.800 ;
        RECT 138.960 165.630 139.310 165.800 ;
        RECT 139.600 165.630 139.950 165.800 ;
        RECT 140.240 165.630 140.590 165.800 ;
        RECT 140.880 165.630 141.230 165.800 ;
        RECT 141.520 165.630 141.870 165.800 ;
        RECT 134.890 159.375 135.060 165.415 ;
        RECT 135.530 159.375 135.700 165.415 ;
        RECT 136.170 159.375 136.340 165.415 ;
        RECT 136.810 159.375 136.980 165.415 ;
        RECT 137.450 159.375 137.620 165.415 ;
        RECT 138.090 159.375 138.260 165.415 ;
        RECT 138.730 159.375 138.900 165.415 ;
        RECT 139.370 159.375 139.540 165.415 ;
        RECT 140.010 159.375 140.180 165.415 ;
        RECT 140.650 159.375 140.820 165.415 ;
        RECT 141.290 159.375 141.460 165.415 ;
        RECT 141.930 159.375 142.100 165.415 ;
        RECT 135.120 158.990 135.470 159.160 ;
        RECT 135.760 158.990 136.110 159.160 ;
        RECT 136.400 158.990 136.750 159.160 ;
        RECT 137.040 158.990 137.390 159.160 ;
        RECT 137.680 158.990 138.030 159.160 ;
        RECT 138.320 158.990 138.670 159.160 ;
        RECT 138.960 158.990 139.310 159.160 ;
        RECT 139.600 158.990 139.950 159.160 ;
        RECT 140.240 158.990 140.590 159.160 ;
        RECT 140.880 158.990 141.230 159.160 ;
        RECT 141.520 158.990 141.870 159.160 ;
        RECT 135.140 158.650 141.090 158.655 ;
        RECT 142.500 158.650 143.390 166.140 ;
        RECT 133.640 158.480 143.390 158.650 ;
        RECT 133.640 156.490 141.090 158.480 ;
        RECT 141.490 157.070 141.660 158.110 ;
        RECT 141.930 157.070 142.100 158.110 ;
        RECT 141.630 156.685 141.960 156.855 ;
        RECT 142.500 156.490 143.390 158.480 ;
        RECT 133.640 155.990 143.390 156.490 ;
        RECT 133.640 148.650 134.490 155.990 ;
        RECT 135.120 155.630 135.470 155.800 ;
        RECT 135.760 155.630 136.110 155.800 ;
        RECT 136.400 155.630 136.750 155.800 ;
        RECT 137.040 155.630 137.390 155.800 ;
        RECT 137.680 155.630 138.030 155.800 ;
        RECT 138.320 155.630 138.670 155.800 ;
        RECT 138.960 155.630 139.310 155.800 ;
        RECT 139.600 155.630 139.950 155.800 ;
        RECT 140.240 155.630 140.590 155.800 ;
        RECT 140.880 155.630 141.230 155.800 ;
        RECT 141.520 155.630 141.870 155.800 ;
        RECT 134.890 149.375 135.060 155.415 ;
        RECT 135.530 149.375 135.700 155.415 ;
        RECT 136.170 149.375 136.340 155.415 ;
        RECT 136.810 149.375 136.980 155.415 ;
        RECT 137.450 149.375 137.620 155.415 ;
        RECT 138.090 149.375 138.260 155.415 ;
        RECT 138.730 149.375 138.900 155.415 ;
        RECT 139.370 149.375 139.540 155.415 ;
        RECT 140.010 149.375 140.180 155.415 ;
        RECT 140.650 149.375 140.820 155.415 ;
        RECT 141.290 149.375 141.460 155.415 ;
        RECT 141.930 149.375 142.100 155.415 ;
        RECT 135.120 148.990 135.470 149.160 ;
        RECT 135.760 148.990 136.110 149.160 ;
        RECT 136.400 148.990 136.750 149.160 ;
        RECT 137.040 148.990 137.390 149.160 ;
        RECT 137.680 148.990 138.030 149.160 ;
        RECT 138.320 148.990 138.670 149.160 ;
        RECT 138.960 148.990 139.310 149.160 ;
        RECT 139.600 148.990 139.950 149.160 ;
        RECT 140.240 148.990 140.590 149.160 ;
        RECT 140.880 148.990 141.230 149.160 ;
        RECT 141.520 148.990 141.870 149.160 ;
        RECT 135.140 148.650 141.090 148.655 ;
        RECT 142.500 148.650 143.390 155.990 ;
        RECT 133.640 148.480 143.390 148.650 ;
        RECT 133.640 146.490 141.090 148.480 ;
        RECT 141.490 147.070 141.660 148.110 ;
        RECT 141.930 147.070 142.100 148.110 ;
        RECT 141.630 146.685 141.960 146.855 ;
        RECT 142.500 146.490 143.390 148.480 ;
        RECT 133.640 145.990 143.390 146.490 ;
        RECT 133.640 138.650 134.490 145.990 ;
        RECT 135.120 145.630 135.470 145.800 ;
        RECT 135.760 145.630 136.110 145.800 ;
        RECT 136.400 145.630 136.750 145.800 ;
        RECT 137.040 145.630 137.390 145.800 ;
        RECT 137.680 145.630 138.030 145.800 ;
        RECT 138.320 145.630 138.670 145.800 ;
        RECT 138.960 145.630 139.310 145.800 ;
        RECT 139.600 145.630 139.950 145.800 ;
        RECT 140.240 145.630 140.590 145.800 ;
        RECT 140.880 145.630 141.230 145.800 ;
        RECT 141.520 145.630 141.870 145.800 ;
        RECT 134.890 139.375 135.060 145.415 ;
        RECT 135.530 139.375 135.700 145.415 ;
        RECT 136.170 139.375 136.340 145.415 ;
        RECT 136.810 139.375 136.980 145.415 ;
        RECT 137.450 139.375 137.620 145.415 ;
        RECT 138.090 139.375 138.260 145.415 ;
        RECT 138.730 139.375 138.900 145.415 ;
        RECT 139.370 139.375 139.540 145.415 ;
        RECT 140.010 139.375 140.180 145.415 ;
        RECT 140.650 139.375 140.820 145.415 ;
        RECT 141.290 139.375 141.460 145.415 ;
        RECT 141.930 139.375 142.100 145.415 ;
        RECT 135.120 138.990 135.470 139.160 ;
        RECT 135.760 138.990 136.110 139.160 ;
        RECT 136.400 138.990 136.750 139.160 ;
        RECT 137.040 138.990 137.390 139.160 ;
        RECT 137.680 138.990 138.030 139.160 ;
        RECT 138.320 138.990 138.670 139.160 ;
        RECT 138.960 138.990 139.310 139.160 ;
        RECT 139.600 138.990 139.950 139.160 ;
        RECT 140.240 138.990 140.590 139.160 ;
        RECT 140.880 138.990 141.230 139.160 ;
        RECT 141.520 138.990 141.870 139.160 ;
        RECT 135.140 138.650 141.090 138.655 ;
        RECT 142.500 138.650 143.390 145.990 ;
        RECT 133.640 138.480 143.390 138.650 ;
        RECT 133.640 136.490 141.090 138.480 ;
        RECT 141.490 137.070 141.660 138.110 ;
        RECT 141.930 137.070 142.100 138.110 ;
        RECT 141.630 136.685 141.960 136.855 ;
        RECT 142.500 136.490 143.390 138.480 ;
        RECT 133.640 135.990 143.390 136.490 ;
        RECT 133.640 128.650 134.490 135.990 ;
        RECT 135.120 135.630 135.470 135.800 ;
        RECT 135.760 135.630 136.110 135.800 ;
        RECT 136.400 135.630 136.750 135.800 ;
        RECT 137.040 135.630 137.390 135.800 ;
        RECT 137.680 135.630 138.030 135.800 ;
        RECT 138.320 135.630 138.670 135.800 ;
        RECT 138.960 135.630 139.310 135.800 ;
        RECT 139.600 135.630 139.950 135.800 ;
        RECT 140.240 135.630 140.590 135.800 ;
        RECT 140.880 135.630 141.230 135.800 ;
        RECT 141.520 135.630 141.870 135.800 ;
        RECT 134.890 129.375 135.060 135.415 ;
        RECT 135.530 129.375 135.700 135.415 ;
        RECT 136.170 129.375 136.340 135.415 ;
        RECT 136.810 129.375 136.980 135.415 ;
        RECT 137.450 129.375 137.620 135.415 ;
        RECT 138.090 129.375 138.260 135.415 ;
        RECT 138.730 129.375 138.900 135.415 ;
        RECT 139.370 129.375 139.540 135.415 ;
        RECT 140.010 129.375 140.180 135.415 ;
        RECT 140.650 129.375 140.820 135.415 ;
        RECT 141.290 129.375 141.460 135.415 ;
        RECT 141.930 129.375 142.100 135.415 ;
        RECT 135.120 128.990 135.470 129.160 ;
        RECT 135.760 128.990 136.110 129.160 ;
        RECT 136.400 128.990 136.750 129.160 ;
        RECT 137.040 128.990 137.390 129.160 ;
        RECT 137.680 128.990 138.030 129.160 ;
        RECT 138.320 128.990 138.670 129.160 ;
        RECT 138.960 128.990 139.310 129.160 ;
        RECT 139.600 128.990 139.950 129.160 ;
        RECT 140.240 128.990 140.590 129.160 ;
        RECT 140.880 128.990 141.230 129.160 ;
        RECT 141.520 128.990 141.870 129.160 ;
        RECT 135.140 128.650 141.090 128.655 ;
        RECT 142.500 128.650 143.390 135.990 ;
        RECT 133.640 128.480 143.390 128.650 ;
        RECT 133.640 126.490 141.090 128.480 ;
        RECT 141.490 127.070 141.660 128.110 ;
        RECT 141.930 127.070 142.100 128.110 ;
        RECT 141.630 126.685 141.960 126.855 ;
        RECT 142.500 126.490 143.390 128.480 ;
        RECT 133.640 125.990 143.390 126.490 ;
        RECT 133.640 118.650 134.490 125.990 ;
        RECT 135.120 125.630 135.470 125.800 ;
        RECT 135.760 125.630 136.110 125.800 ;
        RECT 136.400 125.630 136.750 125.800 ;
        RECT 137.040 125.630 137.390 125.800 ;
        RECT 137.680 125.630 138.030 125.800 ;
        RECT 138.320 125.630 138.670 125.800 ;
        RECT 138.960 125.630 139.310 125.800 ;
        RECT 139.600 125.630 139.950 125.800 ;
        RECT 140.240 125.630 140.590 125.800 ;
        RECT 140.880 125.630 141.230 125.800 ;
        RECT 141.520 125.630 141.870 125.800 ;
        RECT 134.890 119.375 135.060 125.415 ;
        RECT 135.530 119.375 135.700 125.415 ;
        RECT 136.170 119.375 136.340 125.415 ;
        RECT 136.810 119.375 136.980 125.415 ;
        RECT 137.450 119.375 137.620 125.415 ;
        RECT 138.090 119.375 138.260 125.415 ;
        RECT 138.730 119.375 138.900 125.415 ;
        RECT 139.370 119.375 139.540 125.415 ;
        RECT 140.010 119.375 140.180 125.415 ;
        RECT 140.650 119.375 140.820 125.415 ;
        RECT 141.290 119.375 141.460 125.415 ;
        RECT 141.930 119.375 142.100 125.415 ;
        RECT 135.120 118.990 135.470 119.160 ;
        RECT 135.760 118.990 136.110 119.160 ;
        RECT 136.400 118.990 136.750 119.160 ;
        RECT 137.040 118.990 137.390 119.160 ;
        RECT 137.680 118.990 138.030 119.160 ;
        RECT 138.320 118.990 138.670 119.160 ;
        RECT 138.960 118.990 139.310 119.160 ;
        RECT 139.600 118.990 139.950 119.160 ;
        RECT 140.240 118.990 140.590 119.160 ;
        RECT 140.880 118.990 141.230 119.160 ;
        RECT 141.520 118.990 141.870 119.160 ;
        RECT 135.140 118.650 141.090 118.655 ;
        RECT 142.500 118.650 143.390 125.990 ;
        RECT 133.640 118.480 143.390 118.650 ;
        RECT 133.640 116.490 141.090 118.480 ;
        RECT 141.490 117.070 141.660 118.110 ;
        RECT 141.930 117.070 142.100 118.110 ;
        RECT 141.630 116.685 141.960 116.855 ;
        RECT 142.500 116.490 143.390 118.480 ;
        RECT 133.640 115.990 143.390 116.490 ;
        RECT 133.640 108.650 134.490 115.990 ;
        RECT 135.120 115.630 135.470 115.800 ;
        RECT 135.760 115.630 136.110 115.800 ;
        RECT 136.400 115.630 136.750 115.800 ;
        RECT 137.040 115.630 137.390 115.800 ;
        RECT 137.680 115.630 138.030 115.800 ;
        RECT 138.320 115.630 138.670 115.800 ;
        RECT 138.960 115.630 139.310 115.800 ;
        RECT 139.600 115.630 139.950 115.800 ;
        RECT 140.240 115.630 140.590 115.800 ;
        RECT 140.880 115.630 141.230 115.800 ;
        RECT 141.520 115.630 141.870 115.800 ;
        RECT 134.890 109.375 135.060 115.415 ;
        RECT 135.530 109.375 135.700 115.415 ;
        RECT 136.170 109.375 136.340 115.415 ;
        RECT 136.810 109.375 136.980 115.415 ;
        RECT 137.450 109.375 137.620 115.415 ;
        RECT 138.090 109.375 138.260 115.415 ;
        RECT 138.730 109.375 138.900 115.415 ;
        RECT 139.370 109.375 139.540 115.415 ;
        RECT 140.010 109.375 140.180 115.415 ;
        RECT 140.650 109.375 140.820 115.415 ;
        RECT 141.290 109.375 141.460 115.415 ;
        RECT 141.930 109.375 142.100 115.415 ;
        RECT 135.120 108.990 135.470 109.160 ;
        RECT 135.760 108.990 136.110 109.160 ;
        RECT 136.400 108.990 136.750 109.160 ;
        RECT 137.040 108.990 137.390 109.160 ;
        RECT 137.680 108.990 138.030 109.160 ;
        RECT 138.320 108.990 138.670 109.160 ;
        RECT 138.960 108.990 139.310 109.160 ;
        RECT 139.600 108.990 139.950 109.160 ;
        RECT 140.240 108.990 140.590 109.160 ;
        RECT 140.880 108.990 141.230 109.160 ;
        RECT 141.520 108.990 141.870 109.160 ;
        RECT 135.140 108.650 141.090 108.655 ;
        RECT 142.500 108.650 143.390 115.990 ;
        RECT 133.640 108.480 143.390 108.650 ;
        RECT 133.640 106.490 141.090 108.480 ;
        RECT 141.490 107.070 141.660 108.110 ;
        RECT 141.930 107.070 142.100 108.110 ;
        RECT 141.630 106.685 141.960 106.855 ;
        RECT 142.500 106.490 143.390 108.480 ;
        RECT 133.640 105.990 143.390 106.490 ;
        RECT 133.640 98.650 134.490 105.990 ;
        RECT 135.120 105.630 135.470 105.800 ;
        RECT 135.760 105.630 136.110 105.800 ;
        RECT 136.400 105.630 136.750 105.800 ;
        RECT 137.040 105.630 137.390 105.800 ;
        RECT 137.680 105.630 138.030 105.800 ;
        RECT 138.320 105.630 138.670 105.800 ;
        RECT 138.960 105.630 139.310 105.800 ;
        RECT 139.600 105.630 139.950 105.800 ;
        RECT 140.240 105.630 140.590 105.800 ;
        RECT 140.880 105.630 141.230 105.800 ;
        RECT 141.520 105.630 141.870 105.800 ;
        RECT 134.890 99.375 135.060 105.415 ;
        RECT 135.530 99.375 135.700 105.415 ;
        RECT 136.170 99.375 136.340 105.415 ;
        RECT 136.810 99.375 136.980 105.415 ;
        RECT 137.450 99.375 137.620 105.415 ;
        RECT 138.090 99.375 138.260 105.415 ;
        RECT 138.730 99.375 138.900 105.415 ;
        RECT 139.370 99.375 139.540 105.415 ;
        RECT 140.010 99.375 140.180 105.415 ;
        RECT 140.650 99.375 140.820 105.415 ;
        RECT 141.290 99.375 141.460 105.415 ;
        RECT 141.930 99.375 142.100 105.415 ;
        RECT 135.120 98.990 135.470 99.160 ;
        RECT 135.760 98.990 136.110 99.160 ;
        RECT 136.400 98.990 136.750 99.160 ;
        RECT 137.040 98.990 137.390 99.160 ;
        RECT 137.680 98.990 138.030 99.160 ;
        RECT 138.320 98.990 138.670 99.160 ;
        RECT 138.960 98.990 139.310 99.160 ;
        RECT 139.600 98.990 139.950 99.160 ;
        RECT 140.240 98.990 140.590 99.160 ;
        RECT 140.880 98.990 141.230 99.160 ;
        RECT 141.520 98.990 141.870 99.160 ;
        RECT 135.140 98.650 141.090 98.655 ;
        RECT 142.500 98.650 143.390 105.990 ;
        RECT 133.640 98.480 143.390 98.650 ;
        RECT 133.640 96.490 141.090 98.480 ;
        RECT 141.490 97.070 141.660 98.110 ;
        RECT 141.930 97.070 142.100 98.110 ;
        RECT 141.630 96.685 141.960 96.855 ;
        RECT 142.500 96.490 143.390 98.480 ;
        RECT 133.640 95.990 143.390 96.490 ;
        RECT 133.640 88.650 134.490 95.990 ;
        RECT 135.120 95.630 135.470 95.800 ;
        RECT 135.760 95.630 136.110 95.800 ;
        RECT 136.400 95.630 136.750 95.800 ;
        RECT 137.040 95.630 137.390 95.800 ;
        RECT 137.680 95.630 138.030 95.800 ;
        RECT 138.320 95.630 138.670 95.800 ;
        RECT 138.960 95.630 139.310 95.800 ;
        RECT 139.600 95.630 139.950 95.800 ;
        RECT 140.240 95.630 140.590 95.800 ;
        RECT 140.880 95.630 141.230 95.800 ;
        RECT 141.520 95.630 141.870 95.800 ;
        RECT 134.890 89.375 135.060 95.415 ;
        RECT 135.530 89.375 135.700 95.415 ;
        RECT 136.170 89.375 136.340 95.415 ;
        RECT 136.810 89.375 136.980 95.415 ;
        RECT 137.450 89.375 137.620 95.415 ;
        RECT 138.090 89.375 138.260 95.415 ;
        RECT 138.730 89.375 138.900 95.415 ;
        RECT 139.370 89.375 139.540 95.415 ;
        RECT 140.010 89.375 140.180 95.415 ;
        RECT 140.650 89.375 140.820 95.415 ;
        RECT 141.290 89.375 141.460 95.415 ;
        RECT 141.930 89.375 142.100 95.415 ;
        RECT 135.120 88.990 135.470 89.160 ;
        RECT 135.760 88.990 136.110 89.160 ;
        RECT 136.400 88.990 136.750 89.160 ;
        RECT 137.040 88.990 137.390 89.160 ;
        RECT 137.680 88.990 138.030 89.160 ;
        RECT 138.320 88.990 138.670 89.160 ;
        RECT 138.960 88.990 139.310 89.160 ;
        RECT 139.600 88.990 139.950 89.160 ;
        RECT 140.240 88.990 140.590 89.160 ;
        RECT 140.880 88.990 141.230 89.160 ;
        RECT 141.520 88.990 141.870 89.160 ;
        RECT 135.140 88.650 141.090 88.655 ;
        RECT 142.500 88.650 143.390 95.990 ;
        RECT 133.640 88.480 143.390 88.650 ;
        RECT 133.640 86.490 141.090 88.480 ;
        RECT 141.490 87.070 141.660 88.110 ;
        RECT 141.930 87.070 142.100 88.110 ;
        RECT 141.630 86.685 141.960 86.855 ;
        RECT 142.500 86.490 143.390 88.480 ;
        RECT 133.640 85.990 143.390 86.490 ;
        RECT 133.640 78.650 134.490 85.990 ;
        RECT 135.120 85.630 135.470 85.800 ;
        RECT 135.760 85.630 136.110 85.800 ;
        RECT 136.400 85.630 136.750 85.800 ;
        RECT 137.040 85.630 137.390 85.800 ;
        RECT 137.680 85.630 138.030 85.800 ;
        RECT 138.320 85.630 138.670 85.800 ;
        RECT 138.960 85.630 139.310 85.800 ;
        RECT 139.600 85.630 139.950 85.800 ;
        RECT 140.240 85.630 140.590 85.800 ;
        RECT 140.880 85.630 141.230 85.800 ;
        RECT 141.520 85.630 141.870 85.800 ;
        RECT 134.890 79.375 135.060 85.415 ;
        RECT 135.530 79.375 135.700 85.415 ;
        RECT 136.170 79.375 136.340 85.415 ;
        RECT 136.810 79.375 136.980 85.415 ;
        RECT 137.450 79.375 137.620 85.415 ;
        RECT 138.090 79.375 138.260 85.415 ;
        RECT 138.730 79.375 138.900 85.415 ;
        RECT 139.370 79.375 139.540 85.415 ;
        RECT 140.010 79.375 140.180 85.415 ;
        RECT 140.650 79.375 140.820 85.415 ;
        RECT 141.290 79.375 141.460 85.415 ;
        RECT 141.930 79.375 142.100 85.415 ;
        RECT 135.120 78.990 135.470 79.160 ;
        RECT 135.760 78.990 136.110 79.160 ;
        RECT 136.400 78.990 136.750 79.160 ;
        RECT 137.040 78.990 137.390 79.160 ;
        RECT 137.680 78.990 138.030 79.160 ;
        RECT 138.320 78.990 138.670 79.160 ;
        RECT 138.960 78.990 139.310 79.160 ;
        RECT 139.600 78.990 139.950 79.160 ;
        RECT 140.240 78.990 140.590 79.160 ;
        RECT 140.880 78.990 141.230 79.160 ;
        RECT 141.520 78.990 141.870 79.160 ;
        RECT 135.140 78.650 141.090 78.655 ;
        RECT 142.500 78.650 143.390 85.990 ;
        RECT 133.640 78.480 143.390 78.650 ;
        RECT 133.640 76.490 141.090 78.480 ;
        RECT 141.490 77.070 141.660 78.110 ;
        RECT 141.930 77.070 142.100 78.110 ;
        RECT 141.630 76.685 141.960 76.855 ;
        RECT 142.500 76.490 143.390 78.480 ;
        RECT 133.640 75.990 143.390 76.490 ;
        RECT 133.640 68.650 134.490 75.990 ;
        RECT 135.120 75.630 135.470 75.800 ;
        RECT 135.760 75.630 136.110 75.800 ;
        RECT 136.400 75.630 136.750 75.800 ;
        RECT 137.040 75.630 137.390 75.800 ;
        RECT 137.680 75.630 138.030 75.800 ;
        RECT 138.320 75.630 138.670 75.800 ;
        RECT 138.960 75.630 139.310 75.800 ;
        RECT 139.600 75.630 139.950 75.800 ;
        RECT 140.240 75.630 140.590 75.800 ;
        RECT 140.880 75.630 141.230 75.800 ;
        RECT 141.520 75.630 141.870 75.800 ;
        RECT 134.890 69.375 135.060 75.415 ;
        RECT 135.530 69.375 135.700 75.415 ;
        RECT 136.170 69.375 136.340 75.415 ;
        RECT 136.810 69.375 136.980 75.415 ;
        RECT 137.450 69.375 137.620 75.415 ;
        RECT 138.090 69.375 138.260 75.415 ;
        RECT 138.730 69.375 138.900 75.415 ;
        RECT 139.370 69.375 139.540 75.415 ;
        RECT 140.010 69.375 140.180 75.415 ;
        RECT 140.650 69.375 140.820 75.415 ;
        RECT 141.290 69.375 141.460 75.415 ;
        RECT 141.930 69.375 142.100 75.415 ;
        RECT 135.120 68.990 135.470 69.160 ;
        RECT 135.760 68.990 136.110 69.160 ;
        RECT 136.400 68.990 136.750 69.160 ;
        RECT 137.040 68.990 137.390 69.160 ;
        RECT 137.680 68.990 138.030 69.160 ;
        RECT 138.320 68.990 138.670 69.160 ;
        RECT 138.960 68.990 139.310 69.160 ;
        RECT 139.600 68.990 139.950 69.160 ;
        RECT 140.240 68.990 140.590 69.160 ;
        RECT 140.880 68.990 141.230 69.160 ;
        RECT 141.520 68.990 141.870 69.160 ;
        RECT 135.140 68.650 141.090 68.655 ;
        RECT 142.500 68.650 143.390 75.990 ;
        RECT 133.640 68.480 143.390 68.650 ;
        RECT 133.640 66.490 141.090 68.480 ;
        RECT 141.490 67.070 141.660 68.110 ;
        RECT 141.930 67.070 142.100 68.110 ;
        RECT 141.630 66.685 141.960 66.855 ;
        RECT 142.500 66.490 143.390 68.480 ;
        RECT 133.640 65.990 143.390 66.490 ;
        RECT 133.640 58.650 134.490 65.990 ;
        RECT 135.120 65.630 135.470 65.800 ;
        RECT 135.760 65.630 136.110 65.800 ;
        RECT 136.400 65.630 136.750 65.800 ;
        RECT 137.040 65.630 137.390 65.800 ;
        RECT 137.680 65.630 138.030 65.800 ;
        RECT 138.320 65.630 138.670 65.800 ;
        RECT 138.960 65.630 139.310 65.800 ;
        RECT 139.600 65.630 139.950 65.800 ;
        RECT 140.240 65.630 140.590 65.800 ;
        RECT 140.880 65.630 141.230 65.800 ;
        RECT 141.520 65.630 141.870 65.800 ;
        RECT 134.890 59.375 135.060 65.415 ;
        RECT 135.530 59.375 135.700 65.415 ;
        RECT 136.170 59.375 136.340 65.415 ;
        RECT 136.810 59.375 136.980 65.415 ;
        RECT 137.450 59.375 137.620 65.415 ;
        RECT 138.090 59.375 138.260 65.415 ;
        RECT 138.730 59.375 138.900 65.415 ;
        RECT 139.370 59.375 139.540 65.415 ;
        RECT 140.010 59.375 140.180 65.415 ;
        RECT 140.650 59.375 140.820 65.415 ;
        RECT 141.290 59.375 141.460 65.415 ;
        RECT 141.930 59.375 142.100 65.415 ;
        RECT 135.120 58.990 135.470 59.160 ;
        RECT 135.760 58.990 136.110 59.160 ;
        RECT 136.400 58.990 136.750 59.160 ;
        RECT 137.040 58.990 137.390 59.160 ;
        RECT 137.680 58.990 138.030 59.160 ;
        RECT 138.320 58.990 138.670 59.160 ;
        RECT 138.960 58.990 139.310 59.160 ;
        RECT 139.600 58.990 139.950 59.160 ;
        RECT 140.240 58.990 140.590 59.160 ;
        RECT 140.880 58.990 141.230 59.160 ;
        RECT 141.520 58.990 141.870 59.160 ;
        RECT 135.140 58.650 141.090 58.655 ;
        RECT 142.500 58.650 143.390 65.990 ;
        RECT 133.640 58.480 143.390 58.650 ;
        RECT 133.640 56.490 141.090 58.480 ;
        RECT 141.490 57.070 141.660 58.110 ;
        RECT 141.930 57.070 142.100 58.110 ;
        RECT 141.630 56.685 141.960 56.855 ;
        RECT 142.500 56.490 143.390 58.480 ;
        RECT 133.640 55.990 143.390 56.490 ;
        RECT 133.640 48.650 134.490 55.990 ;
        RECT 135.120 55.630 135.470 55.800 ;
        RECT 135.760 55.630 136.110 55.800 ;
        RECT 136.400 55.630 136.750 55.800 ;
        RECT 137.040 55.630 137.390 55.800 ;
        RECT 137.680 55.630 138.030 55.800 ;
        RECT 138.320 55.630 138.670 55.800 ;
        RECT 138.960 55.630 139.310 55.800 ;
        RECT 139.600 55.630 139.950 55.800 ;
        RECT 140.240 55.630 140.590 55.800 ;
        RECT 140.880 55.630 141.230 55.800 ;
        RECT 141.520 55.630 141.870 55.800 ;
        RECT 134.890 49.375 135.060 55.415 ;
        RECT 135.530 49.375 135.700 55.415 ;
        RECT 136.170 49.375 136.340 55.415 ;
        RECT 136.810 49.375 136.980 55.415 ;
        RECT 137.450 49.375 137.620 55.415 ;
        RECT 138.090 49.375 138.260 55.415 ;
        RECT 138.730 49.375 138.900 55.415 ;
        RECT 139.370 49.375 139.540 55.415 ;
        RECT 140.010 49.375 140.180 55.415 ;
        RECT 140.650 49.375 140.820 55.415 ;
        RECT 141.290 49.375 141.460 55.415 ;
        RECT 141.930 49.375 142.100 55.415 ;
        RECT 135.120 48.990 135.470 49.160 ;
        RECT 135.760 48.990 136.110 49.160 ;
        RECT 136.400 48.990 136.750 49.160 ;
        RECT 137.040 48.990 137.390 49.160 ;
        RECT 137.680 48.990 138.030 49.160 ;
        RECT 138.320 48.990 138.670 49.160 ;
        RECT 138.960 48.990 139.310 49.160 ;
        RECT 139.600 48.990 139.950 49.160 ;
        RECT 140.240 48.990 140.590 49.160 ;
        RECT 140.880 48.990 141.230 49.160 ;
        RECT 141.520 48.990 141.870 49.160 ;
        RECT 135.140 48.650 141.090 48.655 ;
        RECT 142.500 48.650 143.390 55.990 ;
        RECT 133.640 48.480 143.390 48.650 ;
        RECT 133.640 46.490 141.090 48.480 ;
        RECT 141.490 47.070 141.660 48.110 ;
        RECT 141.930 47.070 142.100 48.110 ;
        RECT 141.630 46.685 141.960 46.855 ;
        RECT 142.500 46.490 143.390 48.480 ;
        RECT 133.640 45.990 143.390 46.490 ;
        RECT 133.640 38.650 134.490 45.990 ;
        RECT 135.120 45.630 135.470 45.800 ;
        RECT 135.760 45.630 136.110 45.800 ;
        RECT 136.400 45.630 136.750 45.800 ;
        RECT 137.040 45.630 137.390 45.800 ;
        RECT 137.680 45.630 138.030 45.800 ;
        RECT 138.320 45.630 138.670 45.800 ;
        RECT 138.960 45.630 139.310 45.800 ;
        RECT 139.600 45.630 139.950 45.800 ;
        RECT 140.240 45.630 140.590 45.800 ;
        RECT 140.880 45.630 141.230 45.800 ;
        RECT 141.520 45.630 141.870 45.800 ;
        RECT 134.890 39.375 135.060 45.415 ;
        RECT 135.530 39.375 135.700 45.415 ;
        RECT 136.170 39.375 136.340 45.415 ;
        RECT 136.810 39.375 136.980 45.415 ;
        RECT 137.450 39.375 137.620 45.415 ;
        RECT 138.090 39.375 138.260 45.415 ;
        RECT 138.730 39.375 138.900 45.415 ;
        RECT 139.370 39.375 139.540 45.415 ;
        RECT 140.010 39.375 140.180 45.415 ;
        RECT 140.650 39.375 140.820 45.415 ;
        RECT 141.290 39.375 141.460 45.415 ;
        RECT 141.930 39.375 142.100 45.415 ;
        RECT 135.120 38.990 135.470 39.160 ;
        RECT 135.760 38.990 136.110 39.160 ;
        RECT 136.400 38.990 136.750 39.160 ;
        RECT 137.040 38.990 137.390 39.160 ;
        RECT 137.680 38.990 138.030 39.160 ;
        RECT 138.320 38.990 138.670 39.160 ;
        RECT 138.960 38.990 139.310 39.160 ;
        RECT 139.600 38.990 139.950 39.160 ;
        RECT 140.240 38.990 140.590 39.160 ;
        RECT 140.880 38.990 141.230 39.160 ;
        RECT 141.520 38.990 141.870 39.160 ;
        RECT 135.140 38.650 141.090 38.655 ;
        RECT 142.500 38.650 143.390 45.990 ;
        RECT 133.640 38.480 143.390 38.650 ;
        RECT 133.640 36.490 141.090 38.480 ;
        RECT 141.490 37.070 141.660 38.110 ;
        RECT 141.930 37.070 142.100 38.110 ;
        RECT 141.630 36.685 141.960 36.855 ;
        RECT 142.500 36.490 143.390 38.480 ;
        RECT 133.640 35.990 143.390 36.490 ;
        RECT 133.640 28.650 134.490 35.990 ;
        RECT 135.120 35.630 135.470 35.800 ;
        RECT 135.760 35.630 136.110 35.800 ;
        RECT 136.400 35.630 136.750 35.800 ;
        RECT 137.040 35.630 137.390 35.800 ;
        RECT 137.680 35.630 138.030 35.800 ;
        RECT 138.320 35.630 138.670 35.800 ;
        RECT 138.960 35.630 139.310 35.800 ;
        RECT 139.600 35.630 139.950 35.800 ;
        RECT 140.240 35.630 140.590 35.800 ;
        RECT 140.880 35.630 141.230 35.800 ;
        RECT 141.520 35.630 141.870 35.800 ;
        RECT 134.890 29.375 135.060 35.415 ;
        RECT 135.530 29.375 135.700 35.415 ;
        RECT 136.170 29.375 136.340 35.415 ;
        RECT 136.810 29.375 136.980 35.415 ;
        RECT 137.450 29.375 137.620 35.415 ;
        RECT 138.090 29.375 138.260 35.415 ;
        RECT 138.730 29.375 138.900 35.415 ;
        RECT 139.370 29.375 139.540 35.415 ;
        RECT 140.010 29.375 140.180 35.415 ;
        RECT 140.650 29.375 140.820 35.415 ;
        RECT 141.290 29.375 141.460 35.415 ;
        RECT 141.930 29.375 142.100 35.415 ;
        RECT 135.120 28.990 135.470 29.160 ;
        RECT 135.760 28.990 136.110 29.160 ;
        RECT 136.400 28.990 136.750 29.160 ;
        RECT 137.040 28.990 137.390 29.160 ;
        RECT 137.680 28.990 138.030 29.160 ;
        RECT 138.320 28.990 138.670 29.160 ;
        RECT 138.960 28.990 139.310 29.160 ;
        RECT 139.600 28.990 139.950 29.160 ;
        RECT 140.240 28.990 140.590 29.160 ;
        RECT 140.880 28.990 141.230 29.160 ;
        RECT 141.520 28.990 141.870 29.160 ;
        RECT 135.140 28.650 141.090 28.655 ;
        RECT 142.500 28.650 143.390 35.990 ;
        RECT 133.640 28.480 143.390 28.650 ;
        RECT 133.640 26.490 141.090 28.480 ;
        RECT 141.490 27.070 141.660 28.110 ;
        RECT 141.930 27.070 142.100 28.110 ;
        RECT 141.630 26.685 141.960 26.855 ;
        RECT 142.500 26.490 143.390 28.480 ;
        RECT 133.640 25.990 143.390 26.490 ;
        RECT 133.640 18.650 134.490 25.990 ;
        RECT 135.120 25.630 135.470 25.800 ;
        RECT 135.760 25.630 136.110 25.800 ;
        RECT 136.400 25.630 136.750 25.800 ;
        RECT 137.040 25.630 137.390 25.800 ;
        RECT 137.680 25.630 138.030 25.800 ;
        RECT 138.320 25.630 138.670 25.800 ;
        RECT 138.960 25.630 139.310 25.800 ;
        RECT 139.600 25.630 139.950 25.800 ;
        RECT 140.240 25.630 140.590 25.800 ;
        RECT 140.880 25.630 141.230 25.800 ;
        RECT 141.520 25.630 141.870 25.800 ;
        RECT 134.890 19.375 135.060 25.415 ;
        RECT 135.530 19.375 135.700 25.415 ;
        RECT 136.170 19.375 136.340 25.415 ;
        RECT 136.810 19.375 136.980 25.415 ;
        RECT 137.450 19.375 137.620 25.415 ;
        RECT 138.090 19.375 138.260 25.415 ;
        RECT 138.730 19.375 138.900 25.415 ;
        RECT 139.370 19.375 139.540 25.415 ;
        RECT 140.010 19.375 140.180 25.415 ;
        RECT 140.650 19.375 140.820 25.415 ;
        RECT 141.290 19.375 141.460 25.415 ;
        RECT 141.930 19.375 142.100 25.415 ;
        RECT 135.120 18.990 135.470 19.160 ;
        RECT 135.760 18.990 136.110 19.160 ;
        RECT 136.400 18.990 136.750 19.160 ;
        RECT 137.040 18.990 137.390 19.160 ;
        RECT 137.680 18.990 138.030 19.160 ;
        RECT 138.320 18.990 138.670 19.160 ;
        RECT 138.960 18.990 139.310 19.160 ;
        RECT 139.600 18.990 139.950 19.160 ;
        RECT 140.240 18.990 140.590 19.160 ;
        RECT 140.880 18.990 141.230 19.160 ;
        RECT 141.520 18.990 141.870 19.160 ;
        RECT 135.140 18.650 141.090 18.655 ;
        RECT 142.500 18.650 143.390 25.990 ;
        RECT 133.640 18.480 143.390 18.650 ;
        RECT 133.640 16.490 141.090 18.480 ;
        RECT 141.490 17.070 141.660 18.110 ;
        RECT 141.930 17.070 142.100 18.110 ;
        RECT 141.630 16.685 141.960 16.855 ;
        RECT 142.500 16.490 143.390 18.480 ;
        RECT 133.640 15.990 143.390 16.490 ;
        RECT 133.640 8.650 134.490 15.990 ;
        RECT 135.120 15.630 135.470 15.800 ;
        RECT 135.760 15.630 136.110 15.800 ;
        RECT 136.400 15.630 136.750 15.800 ;
        RECT 137.040 15.630 137.390 15.800 ;
        RECT 137.680 15.630 138.030 15.800 ;
        RECT 138.320 15.630 138.670 15.800 ;
        RECT 138.960 15.630 139.310 15.800 ;
        RECT 139.600 15.630 139.950 15.800 ;
        RECT 140.240 15.630 140.590 15.800 ;
        RECT 140.880 15.630 141.230 15.800 ;
        RECT 141.520 15.630 141.870 15.800 ;
        RECT 134.890 9.375 135.060 15.415 ;
        RECT 135.530 9.375 135.700 15.415 ;
        RECT 136.170 9.375 136.340 15.415 ;
        RECT 136.810 9.375 136.980 15.415 ;
        RECT 137.450 9.375 137.620 15.415 ;
        RECT 138.090 9.375 138.260 15.415 ;
        RECT 138.730 9.375 138.900 15.415 ;
        RECT 139.370 9.375 139.540 15.415 ;
        RECT 140.010 9.375 140.180 15.415 ;
        RECT 140.650 9.375 140.820 15.415 ;
        RECT 141.290 9.375 141.460 15.415 ;
        RECT 141.930 9.375 142.100 15.415 ;
        RECT 135.120 8.990 135.470 9.160 ;
        RECT 135.760 8.990 136.110 9.160 ;
        RECT 136.400 8.990 136.750 9.160 ;
        RECT 137.040 8.990 137.390 9.160 ;
        RECT 137.680 8.990 138.030 9.160 ;
        RECT 138.320 8.990 138.670 9.160 ;
        RECT 138.960 8.990 139.310 9.160 ;
        RECT 139.600 8.990 139.950 9.160 ;
        RECT 140.240 8.990 140.590 9.160 ;
        RECT 140.880 8.990 141.230 9.160 ;
        RECT 141.520 8.990 141.870 9.160 ;
        RECT 135.140 8.650 141.090 8.655 ;
        RECT 142.500 8.650 143.390 15.990 ;
        RECT 133.640 8.480 143.390 8.650 ;
        RECT 133.640 6.340 141.090 8.480 ;
        RECT 141.490 7.070 141.660 8.110 ;
        RECT 141.930 7.070 142.100 8.110 ;
        RECT 141.630 6.685 141.960 6.855 ;
        RECT 142.500 6.340 143.390 8.480 ;
        RECT 133.640 5.990 143.390 6.340 ;
        RECT 143.565 164.050 152.005 166.490 ;
        RECT 143.565 158.650 144.450 164.050 ;
        RECT 145.080 163.540 145.430 163.710 ;
        RECT 145.720 163.540 146.070 163.710 ;
        RECT 146.360 163.540 146.710 163.710 ;
        RECT 147.000 163.540 147.350 163.710 ;
        RECT 147.640 163.540 147.990 163.710 ;
        RECT 144.850 159.330 145.020 163.370 ;
        RECT 145.490 159.330 145.660 163.370 ;
        RECT 146.130 159.330 146.300 163.370 ;
        RECT 146.770 159.330 146.940 163.370 ;
        RECT 147.410 159.330 147.580 163.370 ;
        RECT 148.050 159.330 148.220 163.370 ;
        RECT 145.080 158.990 145.430 159.160 ;
        RECT 145.720 158.990 146.070 159.160 ;
        RECT 146.360 158.990 146.710 159.160 ;
        RECT 147.000 158.990 147.350 159.160 ;
        RECT 147.640 158.990 147.990 159.160 ;
        RECT 148.620 158.655 152.005 164.050 ;
        RECT 145.865 158.650 152.005 158.655 ;
        RECT 143.565 158.450 152.005 158.650 ;
        RECT 143.565 156.490 144.450 158.450 ;
        RECT 144.850 157.040 145.020 158.080 ;
        RECT 145.290 157.040 145.460 158.080 ;
        RECT 144.990 156.700 145.320 156.870 ;
        RECT 145.860 156.490 152.005 158.450 ;
        RECT 143.565 154.050 152.005 156.490 ;
        RECT 143.565 148.650 144.450 154.050 ;
        RECT 145.080 153.540 145.430 153.710 ;
        RECT 145.720 153.540 146.070 153.710 ;
        RECT 146.360 153.540 146.710 153.710 ;
        RECT 147.000 153.540 147.350 153.710 ;
        RECT 147.640 153.540 147.990 153.710 ;
        RECT 144.850 149.330 145.020 153.370 ;
        RECT 145.490 149.330 145.660 153.370 ;
        RECT 146.130 149.330 146.300 153.370 ;
        RECT 146.770 149.330 146.940 153.370 ;
        RECT 147.410 149.330 147.580 153.370 ;
        RECT 148.050 149.330 148.220 153.370 ;
        RECT 145.080 148.990 145.430 149.160 ;
        RECT 145.720 148.990 146.070 149.160 ;
        RECT 146.360 148.990 146.710 149.160 ;
        RECT 147.000 148.990 147.350 149.160 ;
        RECT 147.640 148.990 147.990 149.160 ;
        RECT 148.620 148.655 152.005 154.050 ;
        RECT 145.865 148.650 152.005 148.655 ;
        RECT 143.565 148.450 152.005 148.650 ;
        RECT 143.565 146.490 144.450 148.450 ;
        RECT 144.850 147.040 145.020 148.080 ;
        RECT 145.290 147.040 145.460 148.080 ;
        RECT 144.990 146.700 145.320 146.870 ;
        RECT 145.860 146.490 152.005 148.450 ;
        RECT 143.565 144.050 152.005 146.490 ;
        RECT 143.565 138.650 144.450 144.050 ;
        RECT 145.080 143.540 145.430 143.710 ;
        RECT 145.720 143.540 146.070 143.710 ;
        RECT 146.360 143.540 146.710 143.710 ;
        RECT 147.000 143.540 147.350 143.710 ;
        RECT 147.640 143.540 147.990 143.710 ;
        RECT 144.850 139.330 145.020 143.370 ;
        RECT 145.490 139.330 145.660 143.370 ;
        RECT 146.130 139.330 146.300 143.370 ;
        RECT 146.770 139.330 146.940 143.370 ;
        RECT 147.410 139.330 147.580 143.370 ;
        RECT 148.050 139.330 148.220 143.370 ;
        RECT 145.080 138.990 145.430 139.160 ;
        RECT 145.720 138.990 146.070 139.160 ;
        RECT 146.360 138.990 146.710 139.160 ;
        RECT 147.000 138.990 147.350 139.160 ;
        RECT 147.640 138.990 147.990 139.160 ;
        RECT 148.620 138.655 152.005 144.050 ;
        RECT 145.865 138.650 152.005 138.655 ;
        RECT 143.565 138.450 152.005 138.650 ;
        RECT 143.565 136.490 144.450 138.450 ;
        RECT 144.850 137.040 145.020 138.080 ;
        RECT 145.290 137.040 145.460 138.080 ;
        RECT 144.990 136.700 145.320 136.870 ;
        RECT 145.860 136.490 152.005 138.450 ;
        RECT 143.565 134.050 152.005 136.490 ;
        RECT 143.565 128.650 144.450 134.050 ;
        RECT 145.080 133.540 145.430 133.710 ;
        RECT 145.720 133.540 146.070 133.710 ;
        RECT 146.360 133.540 146.710 133.710 ;
        RECT 147.000 133.540 147.350 133.710 ;
        RECT 147.640 133.540 147.990 133.710 ;
        RECT 144.850 129.330 145.020 133.370 ;
        RECT 145.490 129.330 145.660 133.370 ;
        RECT 146.130 129.330 146.300 133.370 ;
        RECT 146.770 129.330 146.940 133.370 ;
        RECT 147.410 129.330 147.580 133.370 ;
        RECT 148.050 129.330 148.220 133.370 ;
        RECT 145.080 128.990 145.430 129.160 ;
        RECT 145.720 128.990 146.070 129.160 ;
        RECT 146.360 128.990 146.710 129.160 ;
        RECT 147.000 128.990 147.350 129.160 ;
        RECT 147.640 128.990 147.990 129.160 ;
        RECT 148.620 128.655 152.005 134.050 ;
        RECT 145.865 128.650 152.005 128.655 ;
        RECT 143.565 128.450 152.005 128.650 ;
        RECT 143.565 126.490 144.450 128.450 ;
        RECT 144.850 127.040 145.020 128.080 ;
        RECT 145.290 127.040 145.460 128.080 ;
        RECT 144.990 126.700 145.320 126.870 ;
        RECT 145.860 126.490 152.005 128.450 ;
        RECT 143.565 124.050 152.005 126.490 ;
        RECT 143.565 118.650 144.450 124.050 ;
        RECT 145.080 123.540 145.430 123.710 ;
        RECT 145.720 123.540 146.070 123.710 ;
        RECT 146.360 123.540 146.710 123.710 ;
        RECT 147.000 123.540 147.350 123.710 ;
        RECT 147.640 123.540 147.990 123.710 ;
        RECT 144.850 119.330 145.020 123.370 ;
        RECT 145.490 119.330 145.660 123.370 ;
        RECT 146.130 119.330 146.300 123.370 ;
        RECT 146.770 119.330 146.940 123.370 ;
        RECT 147.410 119.330 147.580 123.370 ;
        RECT 148.050 119.330 148.220 123.370 ;
        RECT 145.080 118.990 145.430 119.160 ;
        RECT 145.720 118.990 146.070 119.160 ;
        RECT 146.360 118.990 146.710 119.160 ;
        RECT 147.000 118.990 147.350 119.160 ;
        RECT 147.640 118.990 147.990 119.160 ;
        RECT 148.620 118.655 152.005 124.050 ;
        RECT 145.865 118.650 152.005 118.655 ;
        RECT 143.565 118.450 152.005 118.650 ;
        RECT 143.565 116.490 144.450 118.450 ;
        RECT 144.850 117.040 145.020 118.080 ;
        RECT 145.290 117.040 145.460 118.080 ;
        RECT 144.990 116.700 145.320 116.870 ;
        RECT 145.860 116.490 152.005 118.450 ;
        RECT 143.565 114.050 152.005 116.490 ;
        RECT 143.565 108.650 144.450 114.050 ;
        RECT 145.080 113.540 145.430 113.710 ;
        RECT 145.720 113.540 146.070 113.710 ;
        RECT 146.360 113.540 146.710 113.710 ;
        RECT 147.000 113.540 147.350 113.710 ;
        RECT 147.640 113.540 147.990 113.710 ;
        RECT 144.850 109.330 145.020 113.370 ;
        RECT 145.490 109.330 145.660 113.370 ;
        RECT 146.130 109.330 146.300 113.370 ;
        RECT 146.770 109.330 146.940 113.370 ;
        RECT 147.410 109.330 147.580 113.370 ;
        RECT 148.050 109.330 148.220 113.370 ;
        RECT 145.080 108.990 145.430 109.160 ;
        RECT 145.720 108.990 146.070 109.160 ;
        RECT 146.360 108.990 146.710 109.160 ;
        RECT 147.000 108.990 147.350 109.160 ;
        RECT 147.640 108.990 147.990 109.160 ;
        RECT 148.620 108.655 152.005 114.050 ;
        RECT 145.865 108.650 152.005 108.655 ;
        RECT 143.565 108.450 152.005 108.650 ;
        RECT 143.565 106.490 144.450 108.450 ;
        RECT 144.850 107.040 145.020 108.080 ;
        RECT 145.290 107.040 145.460 108.080 ;
        RECT 144.990 106.700 145.320 106.870 ;
        RECT 145.860 106.490 152.005 108.450 ;
        RECT 143.565 104.050 152.005 106.490 ;
        RECT 143.565 98.650 144.450 104.050 ;
        RECT 145.080 103.540 145.430 103.710 ;
        RECT 145.720 103.540 146.070 103.710 ;
        RECT 146.360 103.540 146.710 103.710 ;
        RECT 147.000 103.540 147.350 103.710 ;
        RECT 147.640 103.540 147.990 103.710 ;
        RECT 144.850 99.330 145.020 103.370 ;
        RECT 145.490 99.330 145.660 103.370 ;
        RECT 146.130 99.330 146.300 103.370 ;
        RECT 146.770 99.330 146.940 103.370 ;
        RECT 147.410 99.330 147.580 103.370 ;
        RECT 148.050 99.330 148.220 103.370 ;
        RECT 145.080 98.990 145.430 99.160 ;
        RECT 145.720 98.990 146.070 99.160 ;
        RECT 146.360 98.990 146.710 99.160 ;
        RECT 147.000 98.990 147.350 99.160 ;
        RECT 147.640 98.990 147.990 99.160 ;
        RECT 148.620 98.655 152.005 104.050 ;
        RECT 145.865 98.650 152.005 98.655 ;
        RECT 143.565 98.450 152.005 98.650 ;
        RECT 143.565 96.490 144.450 98.450 ;
        RECT 144.850 97.040 145.020 98.080 ;
        RECT 145.290 97.040 145.460 98.080 ;
        RECT 144.990 96.700 145.320 96.870 ;
        RECT 145.860 96.490 152.005 98.450 ;
        RECT 143.565 94.050 152.005 96.490 ;
        RECT 143.565 88.650 144.450 94.050 ;
        RECT 145.080 93.540 145.430 93.710 ;
        RECT 145.720 93.540 146.070 93.710 ;
        RECT 146.360 93.540 146.710 93.710 ;
        RECT 147.000 93.540 147.350 93.710 ;
        RECT 147.640 93.540 147.990 93.710 ;
        RECT 144.850 89.330 145.020 93.370 ;
        RECT 145.490 89.330 145.660 93.370 ;
        RECT 146.130 89.330 146.300 93.370 ;
        RECT 146.770 89.330 146.940 93.370 ;
        RECT 147.410 89.330 147.580 93.370 ;
        RECT 148.050 89.330 148.220 93.370 ;
        RECT 145.080 88.990 145.430 89.160 ;
        RECT 145.720 88.990 146.070 89.160 ;
        RECT 146.360 88.990 146.710 89.160 ;
        RECT 147.000 88.990 147.350 89.160 ;
        RECT 147.640 88.990 147.990 89.160 ;
        RECT 148.620 88.655 152.005 94.050 ;
        RECT 145.865 88.650 152.005 88.655 ;
        RECT 143.565 88.450 152.005 88.650 ;
        RECT 143.565 86.490 144.450 88.450 ;
        RECT 144.850 87.040 145.020 88.080 ;
        RECT 145.290 87.040 145.460 88.080 ;
        RECT 144.990 86.700 145.320 86.870 ;
        RECT 145.860 86.490 152.005 88.450 ;
        RECT 143.565 84.050 152.005 86.490 ;
        RECT 143.565 78.650 144.450 84.050 ;
        RECT 145.080 83.540 145.430 83.710 ;
        RECT 145.720 83.540 146.070 83.710 ;
        RECT 146.360 83.540 146.710 83.710 ;
        RECT 147.000 83.540 147.350 83.710 ;
        RECT 147.640 83.540 147.990 83.710 ;
        RECT 144.850 79.330 145.020 83.370 ;
        RECT 145.490 79.330 145.660 83.370 ;
        RECT 146.130 79.330 146.300 83.370 ;
        RECT 146.770 79.330 146.940 83.370 ;
        RECT 147.410 79.330 147.580 83.370 ;
        RECT 148.050 79.330 148.220 83.370 ;
        RECT 145.080 78.990 145.430 79.160 ;
        RECT 145.720 78.990 146.070 79.160 ;
        RECT 146.360 78.990 146.710 79.160 ;
        RECT 147.000 78.990 147.350 79.160 ;
        RECT 147.640 78.990 147.990 79.160 ;
        RECT 148.620 78.655 152.005 84.050 ;
        RECT 145.865 78.650 152.005 78.655 ;
        RECT 143.565 78.450 152.005 78.650 ;
        RECT 143.565 76.490 144.450 78.450 ;
        RECT 144.850 77.040 145.020 78.080 ;
        RECT 145.290 77.040 145.460 78.080 ;
        RECT 144.990 76.700 145.320 76.870 ;
        RECT 145.860 76.490 152.005 78.450 ;
        RECT 143.565 74.050 152.005 76.490 ;
        RECT 143.565 68.650 144.450 74.050 ;
        RECT 145.080 73.540 145.430 73.710 ;
        RECT 145.720 73.540 146.070 73.710 ;
        RECT 146.360 73.540 146.710 73.710 ;
        RECT 147.000 73.540 147.350 73.710 ;
        RECT 147.640 73.540 147.990 73.710 ;
        RECT 144.850 69.330 145.020 73.370 ;
        RECT 145.490 69.330 145.660 73.370 ;
        RECT 146.130 69.330 146.300 73.370 ;
        RECT 146.770 69.330 146.940 73.370 ;
        RECT 147.410 69.330 147.580 73.370 ;
        RECT 148.050 69.330 148.220 73.370 ;
        RECT 145.080 68.990 145.430 69.160 ;
        RECT 145.720 68.990 146.070 69.160 ;
        RECT 146.360 68.990 146.710 69.160 ;
        RECT 147.000 68.990 147.350 69.160 ;
        RECT 147.640 68.990 147.990 69.160 ;
        RECT 148.620 68.655 152.005 74.050 ;
        RECT 145.865 68.650 152.005 68.655 ;
        RECT 143.565 68.450 152.005 68.650 ;
        RECT 143.565 66.490 144.450 68.450 ;
        RECT 144.850 67.040 145.020 68.080 ;
        RECT 145.290 67.040 145.460 68.080 ;
        RECT 144.990 66.700 145.320 66.870 ;
        RECT 145.860 66.490 152.005 68.450 ;
        RECT 143.565 64.050 152.005 66.490 ;
        RECT 143.565 58.650 144.450 64.050 ;
        RECT 145.080 63.540 145.430 63.710 ;
        RECT 145.720 63.540 146.070 63.710 ;
        RECT 146.360 63.540 146.710 63.710 ;
        RECT 147.000 63.540 147.350 63.710 ;
        RECT 147.640 63.540 147.990 63.710 ;
        RECT 144.850 59.330 145.020 63.370 ;
        RECT 145.490 59.330 145.660 63.370 ;
        RECT 146.130 59.330 146.300 63.370 ;
        RECT 146.770 59.330 146.940 63.370 ;
        RECT 147.410 59.330 147.580 63.370 ;
        RECT 148.050 59.330 148.220 63.370 ;
        RECT 145.080 58.990 145.430 59.160 ;
        RECT 145.720 58.990 146.070 59.160 ;
        RECT 146.360 58.990 146.710 59.160 ;
        RECT 147.000 58.990 147.350 59.160 ;
        RECT 147.640 58.990 147.990 59.160 ;
        RECT 148.620 58.655 152.005 64.050 ;
        RECT 145.865 58.650 152.005 58.655 ;
        RECT 143.565 58.450 152.005 58.650 ;
        RECT 143.565 56.490 144.450 58.450 ;
        RECT 144.850 57.040 145.020 58.080 ;
        RECT 145.290 57.040 145.460 58.080 ;
        RECT 144.990 56.700 145.320 56.870 ;
        RECT 145.860 56.490 152.005 58.450 ;
        RECT 143.565 54.050 152.005 56.490 ;
        RECT 143.565 48.650 144.450 54.050 ;
        RECT 145.080 53.540 145.430 53.710 ;
        RECT 145.720 53.540 146.070 53.710 ;
        RECT 146.360 53.540 146.710 53.710 ;
        RECT 147.000 53.540 147.350 53.710 ;
        RECT 147.640 53.540 147.990 53.710 ;
        RECT 144.850 49.330 145.020 53.370 ;
        RECT 145.490 49.330 145.660 53.370 ;
        RECT 146.130 49.330 146.300 53.370 ;
        RECT 146.770 49.330 146.940 53.370 ;
        RECT 147.410 49.330 147.580 53.370 ;
        RECT 148.050 49.330 148.220 53.370 ;
        RECT 145.080 48.990 145.430 49.160 ;
        RECT 145.720 48.990 146.070 49.160 ;
        RECT 146.360 48.990 146.710 49.160 ;
        RECT 147.000 48.990 147.350 49.160 ;
        RECT 147.640 48.990 147.990 49.160 ;
        RECT 148.620 48.655 152.005 54.050 ;
        RECT 145.865 48.650 152.005 48.655 ;
        RECT 143.565 48.450 152.005 48.650 ;
        RECT 143.565 46.490 144.450 48.450 ;
        RECT 144.850 47.040 145.020 48.080 ;
        RECT 145.290 47.040 145.460 48.080 ;
        RECT 144.990 46.700 145.320 46.870 ;
        RECT 145.860 46.490 152.005 48.450 ;
        RECT 143.565 44.050 152.005 46.490 ;
        RECT 143.565 38.650 144.450 44.050 ;
        RECT 145.080 43.540 145.430 43.710 ;
        RECT 145.720 43.540 146.070 43.710 ;
        RECT 146.360 43.540 146.710 43.710 ;
        RECT 147.000 43.540 147.350 43.710 ;
        RECT 147.640 43.540 147.990 43.710 ;
        RECT 144.850 39.330 145.020 43.370 ;
        RECT 145.490 39.330 145.660 43.370 ;
        RECT 146.130 39.330 146.300 43.370 ;
        RECT 146.770 39.330 146.940 43.370 ;
        RECT 147.410 39.330 147.580 43.370 ;
        RECT 148.050 39.330 148.220 43.370 ;
        RECT 145.080 38.990 145.430 39.160 ;
        RECT 145.720 38.990 146.070 39.160 ;
        RECT 146.360 38.990 146.710 39.160 ;
        RECT 147.000 38.990 147.350 39.160 ;
        RECT 147.640 38.990 147.990 39.160 ;
        RECT 148.620 38.655 152.005 44.050 ;
        RECT 145.865 38.650 152.005 38.655 ;
        RECT 143.565 38.450 152.005 38.650 ;
        RECT 143.565 36.490 144.450 38.450 ;
        RECT 144.850 37.040 145.020 38.080 ;
        RECT 145.290 37.040 145.460 38.080 ;
        RECT 144.990 36.700 145.320 36.870 ;
        RECT 145.860 36.490 152.005 38.450 ;
        RECT 143.565 34.050 152.005 36.490 ;
        RECT 143.565 28.650 144.450 34.050 ;
        RECT 145.080 33.540 145.430 33.710 ;
        RECT 145.720 33.540 146.070 33.710 ;
        RECT 146.360 33.540 146.710 33.710 ;
        RECT 147.000 33.540 147.350 33.710 ;
        RECT 147.640 33.540 147.990 33.710 ;
        RECT 144.850 29.330 145.020 33.370 ;
        RECT 145.490 29.330 145.660 33.370 ;
        RECT 146.130 29.330 146.300 33.370 ;
        RECT 146.770 29.330 146.940 33.370 ;
        RECT 147.410 29.330 147.580 33.370 ;
        RECT 148.050 29.330 148.220 33.370 ;
        RECT 145.080 28.990 145.430 29.160 ;
        RECT 145.720 28.990 146.070 29.160 ;
        RECT 146.360 28.990 146.710 29.160 ;
        RECT 147.000 28.990 147.350 29.160 ;
        RECT 147.640 28.990 147.990 29.160 ;
        RECT 148.620 28.655 152.005 34.050 ;
        RECT 145.865 28.650 152.005 28.655 ;
        RECT 143.565 28.450 152.005 28.650 ;
        RECT 143.565 26.490 144.450 28.450 ;
        RECT 144.850 27.040 145.020 28.080 ;
        RECT 145.290 27.040 145.460 28.080 ;
        RECT 144.990 26.700 145.320 26.870 ;
        RECT 145.860 26.490 152.005 28.450 ;
        RECT 143.565 24.050 152.005 26.490 ;
        RECT 143.565 18.650 144.450 24.050 ;
        RECT 145.080 23.540 145.430 23.710 ;
        RECT 145.720 23.540 146.070 23.710 ;
        RECT 146.360 23.540 146.710 23.710 ;
        RECT 147.000 23.540 147.350 23.710 ;
        RECT 147.640 23.540 147.990 23.710 ;
        RECT 144.850 19.330 145.020 23.370 ;
        RECT 145.490 19.330 145.660 23.370 ;
        RECT 146.130 19.330 146.300 23.370 ;
        RECT 146.770 19.330 146.940 23.370 ;
        RECT 147.410 19.330 147.580 23.370 ;
        RECT 148.050 19.330 148.220 23.370 ;
        RECT 145.080 18.990 145.430 19.160 ;
        RECT 145.720 18.990 146.070 19.160 ;
        RECT 146.360 18.990 146.710 19.160 ;
        RECT 147.000 18.990 147.350 19.160 ;
        RECT 147.640 18.990 147.990 19.160 ;
        RECT 148.620 18.655 152.005 24.050 ;
        RECT 145.865 18.650 152.005 18.655 ;
        RECT 143.565 18.450 152.005 18.650 ;
        RECT 143.565 16.490 144.450 18.450 ;
        RECT 144.850 17.040 145.020 18.080 ;
        RECT 145.290 17.040 145.460 18.080 ;
        RECT 144.990 16.700 145.320 16.870 ;
        RECT 145.860 16.490 152.005 18.450 ;
        RECT 143.565 14.050 152.005 16.490 ;
        RECT 143.565 8.650 144.450 14.050 ;
        RECT 145.080 13.540 145.430 13.710 ;
        RECT 145.720 13.540 146.070 13.710 ;
        RECT 146.360 13.540 146.710 13.710 ;
        RECT 147.000 13.540 147.350 13.710 ;
        RECT 147.640 13.540 147.990 13.710 ;
        RECT 144.850 9.330 145.020 13.370 ;
        RECT 145.490 9.330 145.660 13.370 ;
        RECT 146.130 9.330 146.300 13.370 ;
        RECT 146.770 9.330 146.940 13.370 ;
        RECT 147.410 9.330 147.580 13.370 ;
        RECT 148.050 9.330 148.220 13.370 ;
        RECT 145.080 8.990 145.430 9.160 ;
        RECT 145.720 8.990 146.070 9.160 ;
        RECT 146.360 8.990 146.710 9.160 ;
        RECT 147.000 8.990 147.350 9.160 ;
        RECT 147.640 8.990 147.990 9.160 ;
        RECT 148.620 8.655 152.005 14.050 ;
        RECT 145.865 8.650 152.005 8.655 ;
        RECT 143.565 8.450 152.005 8.650 ;
        RECT 143.565 6.360 144.450 8.450 ;
        RECT 144.850 7.040 145.020 8.080 ;
        RECT 145.290 7.040 145.460 8.080 ;
        RECT 144.990 6.700 145.320 6.870 ;
        RECT 145.860 6.360 152.005 8.450 ;
        RECT 143.565 5.990 152.005 6.360 ;
      LAYER met1 ;
        RECT 78.730 223.870 79.050 223.930 ;
        RECT 116.450 223.870 116.770 223.930 ;
        RECT 78.730 223.730 116.770 223.870 ;
        RECT 78.730 223.670 79.050 223.730 ;
        RECT 116.450 223.670 116.770 223.730 ;
        RECT 117.370 223.870 117.690 223.930 ;
        RECT 151.870 223.870 152.190 223.930 ;
        RECT 117.370 223.730 152.190 223.870 ;
        RECT 117.370 223.670 117.690 223.730 ;
        RECT 151.870 223.670 152.190 223.730 ;
        RECT 2.760 222.800 159.040 223.280 ;
        RECT 4.210 222.310 4.530 222.570 ;
        RECT 7.890 222.310 8.210 222.570 ;
        RECT 11.570 222.310 11.890 222.570 ;
        RECT 16.170 222.310 16.490 222.570 ;
        RECT 18.930 222.310 19.250 222.570 ;
        RECT 22.610 222.310 22.930 222.570 ;
        RECT 26.290 222.310 26.610 222.570 ;
        RECT 29.970 222.310 30.290 222.570 ;
        RECT 69.530 222.510 69.850 222.570 ;
        RECT 59.500 222.370 70.220 222.510 ;
        RECT 48.370 222.170 48.690 222.230 ;
        RECT 58.045 222.170 58.335 222.215 ;
        RECT 48.370 222.030 58.335 222.170 ;
        RECT 48.370 221.970 48.690 222.030 ;
        RECT 58.045 221.985 58.335 222.030 ;
        RECT 59.500 221.980 59.640 222.370 ;
        RECT 69.530 222.310 69.850 222.370 ;
        RECT 64.485 222.170 64.775 222.215 ;
        RECT 66.770 222.170 67.090 222.230 ;
        RECT 64.485 222.030 67.090 222.170 ;
        RECT 70.080 222.170 70.220 222.370 ;
        RECT 70.450 222.310 70.770 222.570 ;
        RECT 77.825 222.510 78.115 222.555 ;
        RECT 78.270 222.510 78.590 222.570 ;
        RECT 89.310 222.510 89.630 222.570 ;
        RECT 77.825 222.370 78.590 222.510 ;
        RECT 77.825 222.325 78.115 222.370 ;
        RECT 78.270 222.310 78.590 222.370 ;
        RECT 82.960 222.370 89.630 222.510 ;
        RECT 71.830 222.170 72.150 222.230 ;
        RECT 70.080 222.030 72.150 222.170 ;
        RECT 59.425 221.750 59.715 221.980 ;
        RECT 61.725 221.935 62.015 221.980 ;
        RECT 63.090 221.935 63.410 221.995 ;
        RECT 64.485 221.985 64.775 222.030 ;
        RECT 66.770 221.970 67.090 222.030 ;
        RECT 71.830 221.970 72.150 222.030 ;
        RECT 61.725 221.795 63.410 221.935 ;
        RECT 61.725 221.750 62.015 221.795 ;
        RECT 63.090 221.735 63.410 221.795 ;
        RECT 65.865 221.830 66.155 221.875 ;
        RECT 67.690 221.830 68.010 221.890 ;
        RECT 65.865 221.690 68.010 221.830 ;
        RECT 68.395 221.725 68.685 221.955 ;
        RECT 65.865 221.645 66.155 221.690 ;
        RECT 67.690 221.630 68.010 221.690 ;
        RECT 63.440 221.490 63.730 221.535 ;
        RECT 64.025 221.490 64.315 221.535 ;
        RECT 66.310 221.490 66.630 221.550 ;
        RECT 63.440 221.305 63.780 221.490 ;
        RECT 64.025 221.350 66.630 221.490 ;
        RECT 64.025 221.305 64.315 221.350 ;
        RECT 62.630 220.950 62.950 221.210 ;
        RECT 63.640 221.150 63.780 221.305 ;
        RECT 66.310 221.290 66.630 221.350 ;
        RECT 66.770 221.490 67.090 221.550 ;
        RECT 68.470 221.490 68.610 221.725 ;
        RECT 69.070 221.710 69.390 221.970 ;
        RECT 77.365 221.950 77.655 221.995 ;
        RECT 77.810 221.950 78.130 222.010 ;
        RECT 71.370 221.630 71.690 221.890 ;
        RECT 77.365 221.810 78.130 221.950 ;
        RECT 77.365 221.765 77.655 221.810 ;
        RECT 77.810 221.750 78.130 221.810 ;
        RECT 78.730 221.800 79.050 222.060 ;
        RECT 81.490 221.935 81.810 221.995 ;
        RECT 82.425 221.935 82.715 221.980 ;
        RECT 82.960 221.935 83.100 222.370 ;
        RECT 89.310 222.310 89.630 222.370 ;
        RECT 90.245 222.510 90.535 222.555 ;
        RECT 95.305 222.510 95.595 222.555 ;
        RECT 90.245 222.370 95.595 222.510 ;
        RECT 90.245 222.325 90.535 222.370 ;
        RECT 95.305 222.325 95.595 222.370 ;
        RECT 95.750 222.510 96.070 222.570 ;
        RECT 98.050 222.510 98.370 222.570 ;
        RECT 116.925 222.510 117.215 222.555 ;
        RECT 136.705 222.510 136.995 222.555 ;
        RECT 142.225 222.510 142.515 222.555 ;
        RECT 155.550 222.510 155.870 222.570 ;
        RECT 95.750 222.370 97.820 222.510 ;
        RECT 95.750 222.310 96.070 222.370 ;
        RECT 81.490 221.795 83.100 221.935 ;
        RECT 81.490 221.735 81.810 221.795 ;
        RECT 82.425 221.750 82.715 221.795 ;
        RECT 84.250 221.735 84.570 221.995 ;
        RECT 85.170 221.970 85.490 222.230 ;
        RECT 97.680 222.170 97.820 222.370 ;
        RECT 98.050 222.370 117.215 222.510 ;
        RECT 98.050 222.310 98.370 222.370 ;
        RECT 116.925 222.325 117.215 222.370 ;
        RECT 124.360 222.370 136.460 222.510 ;
        RECT 109.090 222.170 109.410 222.230 ;
        RECT 124.360 222.170 124.500 222.370 ;
        RECT 86.090 221.830 86.410 221.890 ;
        RECT 87.025 221.830 87.315 221.875 ;
        RECT 86.090 221.690 87.315 221.830 ;
        RECT 94.385 221.830 94.675 222.045 ;
        RECT 97.680 222.030 109.410 222.170 ;
        RECT 109.090 221.970 109.410 222.030 ;
        RECT 115.620 222.030 124.500 222.170 ;
        RECT 124.745 222.170 125.035 222.215 ;
        RECT 132.550 222.170 132.870 222.230 ;
        RECT 124.745 222.030 132.870 222.170 ;
        RECT 136.320 222.170 136.460 222.370 ;
        RECT 136.705 222.370 142.515 222.510 ;
        RECT 136.705 222.325 136.995 222.370 ;
        RECT 142.225 222.325 142.515 222.370 ;
        RECT 146.440 222.370 155.870 222.510 ;
        RECT 146.440 222.170 146.580 222.370 ;
        RECT 155.550 222.310 155.870 222.370 ;
        RECT 136.320 222.030 146.580 222.170 ;
        RECT 146.825 222.170 147.115 222.215 ;
        RECT 153.265 222.170 153.555 222.215 ;
        RECT 146.825 222.030 153.555 222.170 ;
        RECT 94.830 221.830 95.150 221.890 ;
        RECT 94.385 221.815 95.150 221.830 ;
        RECT 94.460 221.690 95.150 221.815 ;
        RECT 86.090 221.630 86.410 221.690 ;
        RECT 87.025 221.645 87.315 221.690 ;
        RECT 94.830 221.630 95.150 221.690 ;
        RECT 95.290 221.870 95.610 221.930 ;
        RECT 95.765 221.870 96.055 221.915 ;
        RECT 95.290 221.730 96.055 221.870 ;
        RECT 95.290 221.670 95.610 221.730 ;
        RECT 95.765 221.685 96.055 221.730 ;
        RECT 96.210 221.670 96.530 221.930 ;
        RECT 109.550 221.630 109.870 221.890 ;
        RECT 110.025 221.685 110.315 221.915 ;
        RECT 110.470 221.830 110.790 221.890 ;
        RECT 113.705 221.830 113.995 221.875 ;
        RECT 115.070 221.830 115.390 221.890 ;
        RECT 115.620 221.875 115.760 222.030 ;
        RECT 124.745 221.985 125.035 222.030 ;
        RECT 132.550 221.970 132.870 222.030 ;
        RECT 146.825 221.985 147.115 222.030 ;
        RECT 153.265 221.985 153.555 222.030 ;
        RECT 110.470 221.690 115.390 221.830 ;
        RECT 74.590 221.490 74.910 221.550 ;
        RECT 66.770 221.350 74.910 221.490 ;
        RECT 66.770 221.290 67.090 221.350 ;
        RECT 74.590 221.290 74.910 221.350 ;
        RECT 77.350 221.490 77.670 221.550 ;
        RECT 108.630 221.490 108.950 221.550 ;
        RECT 77.350 221.350 108.950 221.490 ;
        RECT 77.350 221.290 77.670 221.350 ;
        RECT 108.630 221.290 108.950 221.350 ;
        RECT 110.100 221.210 110.240 221.685 ;
        RECT 110.470 221.630 110.790 221.690 ;
        RECT 113.705 221.645 113.995 221.690 ;
        RECT 115.070 221.630 115.390 221.690 ;
        RECT 115.545 221.645 115.835 221.875 ;
        RECT 115.990 221.630 116.310 221.890 ;
        RECT 123.825 221.645 124.115 221.875 ;
        RECT 120.590 221.490 120.910 221.550 ;
        RECT 122.905 221.490 123.195 221.535 ;
        RECT 120.590 221.350 123.195 221.490 ;
        RECT 123.900 221.490 124.040 221.645 ;
        RECT 126.110 221.630 126.430 221.890 ;
        RECT 127.490 221.630 127.810 221.890 ;
        RECT 133.930 221.630 134.250 221.890 ;
        RECT 136.245 221.830 136.535 221.875 ;
        RECT 138.545 221.830 138.835 221.875 ;
        RECT 136.245 221.690 138.835 221.830 ;
        RECT 136.245 221.645 136.535 221.690 ;
        RECT 138.545 221.645 138.835 221.690 ;
        RECT 139.910 221.830 140.230 221.890 ;
        RECT 141.305 221.830 141.595 221.875 ;
        RECT 139.910 221.690 141.595 221.830 ;
        RECT 139.910 221.630 140.230 221.690 ;
        RECT 141.305 221.645 141.595 221.690 ;
        RECT 143.130 221.630 143.450 221.890 ;
        RECT 150.965 221.830 151.255 221.875 ;
        RECT 152.330 221.830 152.650 221.890 ;
        RECT 145.520 221.690 149.800 221.830 ;
        RECT 126.585 221.490 126.875 221.535 ;
        RECT 123.900 221.350 126.875 221.490 ;
        RECT 120.590 221.290 120.910 221.350 ;
        RECT 122.905 221.305 123.195 221.350 ;
        RECT 126.585 221.305 126.875 221.350 ;
        RECT 131.170 221.490 131.490 221.550 ;
        RECT 137.165 221.490 137.455 221.535 ;
        RECT 137.610 221.490 137.930 221.550 ;
        RECT 145.520 221.535 145.660 221.690 ;
        RECT 145.445 221.490 145.735 221.535 ;
        RECT 131.170 221.350 145.735 221.490 ;
        RECT 65.850 221.150 66.170 221.210 ;
        RECT 63.640 221.010 66.170 221.150 ;
        RECT 65.850 220.950 66.170 221.010 ;
        RECT 69.070 220.950 69.390 221.210 ;
        RECT 79.665 221.150 79.955 221.195 ;
        RECT 81.950 221.150 82.270 221.210 ;
        RECT 79.665 221.010 82.270 221.150 ;
        RECT 79.665 220.965 79.955 221.010 ;
        RECT 81.950 220.950 82.270 221.010 ;
        RECT 82.870 221.150 83.190 221.210 ;
        RECT 93.465 221.150 93.755 221.195 ;
        RECT 82.870 221.010 93.755 221.150 ;
        RECT 82.870 220.950 83.190 221.010 ;
        RECT 93.465 220.965 93.755 221.010 ;
        RECT 96.670 220.950 96.990 221.210 ;
        RECT 106.345 221.150 106.635 221.195 ;
        RECT 108.170 221.150 108.490 221.210 ;
        RECT 106.345 221.010 108.490 221.150 ;
        RECT 106.345 220.965 106.635 221.010 ;
        RECT 108.170 220.950 108.490 221.010 ;
        RECT 110.010 220.950 110.330 221.210 ;
        RECT 110.470 220.950 110.790 221.210 ;
        RECT 122.980 221.150 123.120 221.305 ;
        RECT 131.170 221.290 131.490 221.350 ;
        RECT 137.165 221.305 137.455 221.350 ;
        RECT 137.610 221.290 137.930 221.350 ;
        RECT 145.445 221.305 145.735 221.350 ;
        RECT 145.890 221.490 146.210 221.550 ;
        RECT 149.660 221.535 149.800 221.690 ;
        RECT 150.965 221.690 152.650 221.830 ;
        RECT 150.965 221.645 151.255 221.690 ;
        RECT 152.330 221.630 152.650 221.690 ;
        RECT 152.790 221.830 153.110 221.890 ;
        RECT 156.025 221.830 156.315 221.875 ;
        RECT 152.790 221.690 156.315 221.830 ;
        RECT 152.790 221.630 153.110 221.690 ;
        RECT 156.025 221.645 156.315 221.690 ;
        RECT 146.365 221.490 146.655 221.535 ;
        RECT 145.890 221.350 146.655 221.490 ;
        RECT 145.890 221.290 146.210 221.350 ;
        RECT 146.365 221.305 146.655 221.350 ;
        RECT 149.585 221.305 149.875 221.535 ;
        RECT 150.505 221.490 150.795 221.535 ;
        RECT 154.170 221.490 154.490 221.550 ;
        RECT 150.505 221.350 154.490 221.490 ;
        RECT 150.505 221.305 150.795 221.350 ;
        RECT 154.170 221.290 154.490 221.350 ;
        RECT 125.205 221.150 125.495 221.195 ;
        RECT 122.980 221.010 125.495 221.150 ;
        RECT 125.205 220.965 125.495 221.010 ;
        RECT 133.010 220.950 133.330 221.210 ;
        RECT 134.405 221.150 134.695 221.195 ;
        RECT 135.310 221.150 135.630 221.210 ;
        RECT 134.405 221.010 135.630 221.150 ;
        RECT 134.405 220.965 134.695 221.010 ;
        RECT 135.310 220.950 135.630 221.010 ;
        RECT 147.270 221.150 147.590 221.210 ;
        RECT 148.665 221.150 148.955 221.195 ;
        RECT 147.270 221.010 148.955 221.150 ;
        RECT 147.270 220.950 147.590 221.010 ;
        RECT 148.665 220.965 148.955 221.010 ;
        RECT 152.790 220.950 153.110 221.210 ;
        RECT 1.000 220.080 158.240 220.560 ;
        RECT 76.445 219.790 76.735 219.835 ;
        RECT 64.560 219.650 76.735 219.790 ;
        RECT 58.990 219.540 59.280 219.585 ;
        RECT 61.090 219.540 61.380 219.585 ;
        RECT 62.660 219.540 62.950 219.585 ;
        RECT 58.990 219.400 62.950 219.540 ;
        RECT 58.990 219.355 59.280 219.400 ;
        RECT 61.090 219.355 61.380 219.400 ;
        RECT 62.660 219.355 62.950 219.400 ;
        RECT 59.385 219.200 59.675 219.245 ;
        RECT 60.575 219.200 60.865 219.245 ;
        RECT 63.095 219.200 63.385 219.245 ;
        RECT 54.825 219.110 55.115 219.155 ;
        RECT 58.505 219.110 58.795 219.155 ;
        RECT 54.825 218.970 58.795 219.110 ;
        RECT 59.385 219.060 63.385 219.200 ;
        RECT 59.385 219.015 59.675 219.060 ;
        RECT 60.575 219.015 60.865 219.060 ;
        RECT 63.095 219.015 63.385 219.060 ;
        RECT 54.825 218.925 55.115 218.970 ;
        RECT 58.505 218.925 58.795 218.970 ;
        RECT 54.365 218.770 54.655 218.875 ;
        RECT 56.650 218.770 56.970 218.830 ;
        RECT 54.365 218.645 56.970 218.770 ;
        RECT 54.440 218.630 56.970 218.645 ;
        RECT 56.650 218.570 56.970 218.630 ;
        RECT 57.570 218.570 57.890 218.830 ;
        RECT 59.840 218.770 60.130 218.815 ;
        RECT 64.560 218.770 64.700 219.650 ;
        RECT 76.445 219.605 76.735 219.650 ;
        RECT 86.090 219.590 86.410 219.850 ;
        RECT 107.265 219.790 107.555 219.835 ;
        RECT 110.010 219.790 110.330 219.850 ;
        RECT 107.265 219.650 110.330 219.790 ;
        RECT 107.265 219.605 107.555 219.650 ;
        RECT 110.010 219.590 110.330 219.650 ;
        RECT 118.290 219.590 118.610 219.850 ;
        RECT 137.610 219.790 137.930 219.850 ;
        RECT 140.370 219.790 140.690 219.850 ;
        RECT 144.510 219.790 144.830 219.850 ;
        RECT 137.610 219.650 140.140 219.790 ;
        RECT 137.610 219.590 137.930 219.650 ;
        RECT 79.690 219.540 79.980 219.585 ;
        RECT 81.790 219.540 82.080 219.585 ;
        RECT 83.360 219.540 83.650 219.585 ;
        RECT 59.840 218.630 64.700 218.770 ;
        RECT 65.020 219.310 75.240 219.450 ;
        RECT 79.690 219.400 83.650 219.540 ;
        RECT 100.850 219.540 101.140 219.585 ;
        RECT 102.950 219.540 103.240 219.585 ;
        RECT 104.520 219.540 104.810 219.585 ;
        RECT 95.290 219.450 95.610 219.510 ;
        RECT 99.430 219.450 99.750 219.510 ;
        RECT 79.690 219.355 79.980 219.400 ;
        RECT 81.790 219.355 82.080 219.400 ;
        RECT 83.360 219.355 83.650 219.400 ;
        RECT 59.840 218.585 60.130 218.630 ;
        RECT 56.190 218.230 56.510 218.490 ;
        RECT 56.740 218.430 56.880 218.570 ;
        RECT 65.020 218.430 65.160 219.310 ;
        RECT 67.705 219.110 67.995 219.155 ;
        RECT 69.990 219.110 70.310 219.170 ;
        RECT 67.705 218.970 70.310 219.110 ;
        RECT 67.705 218.925 67.995 218.970 ;
        RECT 69.990 218.910 70.310 218.970 ;
        RECT 75.100 218.955 75.240 219.310 ;
        RECT 84.315 219.310 99.750 219.450 ;
        RECT 100.850 219.400 104.810 219.540 ;
        RECT 110.470 219.540 110.760 219.585 ;
        RECT 112.040 219.540 112.330 219.585 ;
        RECT 114.140 219.540 114.430 219.585 ;
        RECT 100.850 219.355 101.140 219.400 ;
        RECT 102.950 219.355 103.240 219.400 ;
        RECT 104.520 219.355 104.810 219.400 ;
        RECT 107.725 219.450 108.015 219.495 ;
        RECT 109.550 219.450 109.870 219.510 ;
        RECT 80.085 219.200 80.375 219.245 ;
        RECT 81.275 219.200 81.565 219.245 ;
        RECT 83.795 219.200 84.085 219.245 ;
        RECT 75.525 219.110 75.815 219.155 ;
        RECT 79.205 219.110 79.495 219.155 ;
        RECT 75.525 218.970 79.495 219.110 ;
        RECT 80.085 219.060 84.085 219.200 ;
        RECT 80.085 219.015 80.375 219.060 ;
        RECT 81.275 219.015 81.565 219.060 ;
        RECT 83.795 219.015 84.085 219.060 ;
        RECT 69.545 218.770 69.835 218.815 ;
        RECT 70.910 218.770 71.230 218.830 ;
        RECT 69.545 218.630 71.230 218.770 ;
        RECT 71.830 218.645 72.150 218.905 ;
        RECT 74.145 218.660 74.435 218.890 ;
        RECT 75.025 218.770 75.315 218.955 ;
        RECT 75.525 218.925 75.815 218.970 ;
        RECT 79.205 218.925 79.495 218.970 ;
        RECT 76.890 218.770 77.210 218.830 ;
        RECT 75.025 218.725 77.210 218.770 ;
        RECT 69.545 218.585 69.835 218.630 ;
        RECT 70.910 218.570 71.230 218.630 ;
        RECT 56.740 218.290 65.160 218.430 ;
        RECT 65.405 218.430 65.695 218.475 ;
        RECT 65.850 218.430 66.170 218.490 ;
        RECT 65.405 218.290 66.170 218.430 ;
        RECT 65.405 218.245 65.695 218.290 ;
        RECT 65.850 218.230 66.170 218.290 ;
        RECT 69.990 218.430 70.310 218.490 ;
        RECT 72.290 218.430 72.610 218.490 ;
        RECT 69.990 218.290 72.610 218.430 ;
        RECT 69.990 218.230 70.310 218.290 ;
        RECT 72.290 218.230 72.610 218.290 ;
        RECT 73.670 218.230 73.990 218.490 ;
        RECT 74.220 218.430 74.360 218.660 ;
        RECT 75.100 218.630 77.210 218.725 ;
        RECT 76.890 218.570 77.210 218.630 ;
        RECT 77.350 218.570 77.670 218.830 ;
        RECT 77.810 218.770 78.130 218.830 ;
        RECT 78.745 218.770 79.035 218.815 ;
        RECT 77.810 218.630 79.035 218.770 ;
        RECT 77.810 218.570 78.130 218.630 ;
        RECT 78.745 218.585 79.035 218.630 ;
        RECT 80.540 218.770 80.830 218.815 ;
        RECT 82.870 218.770 83.190 218.830 ;
        RECT 80.540 218.630 83.190 218.770 ;
        RECT 80.540 218.585 80.830 218.630 ;
        RECT 75.970 218.430 76.290 218.490 ;
        RECT 74.220 218.290 76.290 218.430 ;
        RECT 75.970 218.230 76.290 218.290 ;
        RECT 76.430 218.430 76.750 218.490 ;
        RECT 78.285 218.430 78.575 218.475 ;
        RECT 76.430 218.290 78.575 218.430 ;
        RECT 78.820 218.430 78.960 218.585 ;
        RECT 82.870 218.570 83.190 218.630 ;
        RECT 84.315 218.430 84.455 219.310 ;
        RECT 95.290 219.250 95.610 219.310 ;
        RECT 99.430 219.250 99.750 219.310 ;
        RECT 107.725 219.310 109.870 219.450 ;
        RECT 110.470 219.400 114.430 219.540 ;
        RECT 122.010 219.540 122.300 219.585 ;
        RECT 124.110 219.540 124.400 219.585 ;
        RECT 125.680 219.540 125.970 219.585 ;
        RECT 110.470 219.355 110.760 219.400 ;
        RECT 112.040 219.355 112.330 219.400 ;
        RECT 114.140 219.355 114.430 219.400 ;
        RECT 115.990 219.450 116.310 219.510 ;
        RECT 107.725 219.265 108.015 219.310 ;
        RECT 109.550 219.250 109.870 219.310 ;
        RECT 115.990 219.310 121.740 219.450 ;
        RECT 122.010 219.400 125.970 219.540 ;
        RECT 122.010 219.355 122.300 219.400 ;
        RECT 124.110 219.355 124.400 219.400 ;
        RECT 125.680 219.355 125.970 219.400 ;
        RECT 133.510 219.540 133.800 219.585 ;
        RECT 135.610 219.540 135.900 219.585 ;
        RECT 137.180 219.540 137.470 219.585 ;
        RECT 133.510 219.400 137.470 219.540 ;
        RECT 133.510 219.355 133.800 219.400 ;
        RECT 135.610 219.355 135.900 219.400 ;
        RECT 137.180 219.355 137.470 219.400 ;
        RECT 140.000 219.450 140.140 219.650 ;
        RECT 140.370 219.650 144.830 219.790 ;
        RECT 140.370 219.590 140.690 219.650 ;
        RECT 144.510 219.590 144.830 219.650 ;
        RECT 151.870 219.590 152.190 219.850 ;
        RECT 152.330 219.790 152.650 219.850 ;
        RECT 152.805 219.790 153.095 219.835 ;
        RECT 152.330 219.650 153.095 219.790 ;
        RECT 152.330 219.590 152.650 219.650 ;
        RECT 152.805 219.605 153.095 219.650 ;
        RECT 145.470 219.540 145.760 219.585 ;
        RECT 147.570 219.540 147.860 219.585 ;
        RECT 149.140 219.540 149.430 219.585 ;
        RECT 140.000 219.310 141.060 219.450 ;
        RECT 145.470 219.400 149.430 219.540 ;
        RECT 145.470 219.355 145.760 219.400 ;
        RECT 147.570 219.355 147.860 219.400 ;
        RECT 149.140 219.355 149.430 219.400 ;
        RECT 115.990 219.250 116.310 219.310 ;
        RECT 101.245 219.200 101.535 219.245 ;
        RECT 102.435 219.200 102.725 219.245 ;
        RECT 104.955 219.200 105.245 219.245 ;
        RECT 87.010 218.910 87.330 219.170 ;
        RECT 89.770 219.110 90.090 219.170 ;
        RECT 93.465 219.110 93.755 219.155 ;
        RECT 89.770 218.970 93.755 219.110 ;
        RECT 89.770 218.910 90.090 218.970 ;
        RECT 93.465 218.925 93.755 218.970 ;
        RECT 98.510 219.110 98.830 219.170 ;
        RECT 98.510 218.970 100.580 219.110 ;
        RECT 101.245 219.060 105.245 219.200 ;
        RECT 110.035 219.200 110.325 219.245 ;
        RECT 112.555 219.200 112.845 219.245 ;
        RECT 113.745 219.200 114.035 219.245 ;
        RECT 108.170 219.110 108.490 219.170 ;
        RECT 101.245 219.015 101.535 219.060 ;
        RECT 102.435 219.015 102.725 219.060 ;
        RECT 104.955 219.015 105.245 219.060 ;
        RECT 98.510 218.910 98.830 218.970 ;
        RECT 87.930 218.645 88.250 218.905 ;
        RECT 89.310 218.645 89.630 218.905 ;
        RECT 96.685 218.770 96.975 218.815 ;
        RECT 96.685 218.630 97.820 218.770 ;
        RECT 96.685 218.585 96.975 218.630 ;
        RECT 78.820 218.290 84.455 218.430 ;
        RECT 93.910 218.430 94.230 218.490 ;
        RECT 97.145 218.430 97.435 218.475 ;
        RECT 93.910 218.290 97.435 218.430 ;
        RECT 97.680 218.430 97.820 218.630 ;
        RECT 98.050 218.570 98.370 218.830 ;
        RECT 99.430 218.570 99.750 218.830 ;
        RECT 100.440 218.815 100.580 218.970 ;
        RECT 105.500 218.970 108.490 219.110 ;
        RECT 110.035 219.060 114.035 219.200 ;
        RECT 110.035 219.015 110.325 219.060 ;
        RECT 112.555 219.015 112.845 219.060 ;
        RECT 113.745 219.015 114.035 219.060 ;
        RECT 114.610 219.110 114.930 219.170 ;
        RECT 121.600 219.110 121.740 219.310 ;
        RECT 122.405 219.200 122.695 219.245 ;
        RECT 123.595 219.200 123.885 219.245 ;
        RECT 126.115 219.200 126.405 219.245 ;
        RECT 100.365 218.585 100.655 218.815 ;
        RECT 101.700 218.770 101.990 218.815 ;
        RECT 105.500 218.770 105.640 218.970 ;
        RECT 108.170 218.910 108.490 218.970 ;
        RECT 114.610 218.970 119.900 219.110 ;
        RECT 121.600 218.970 122.200 219.110 ;
        RECT 122.405 219.060 126.405 219.200 ;
        RECT 122.405 219.015 122.695 219.060 ;
        RECT 123.595 219.015 123.885 219.060 ;
        RECT 126.115 219.015 126.405 219.060 ;
        RECT 133.905 219.200 134.195 219.245 ;
        RECT 135.095 219.200 135.385 219.245 ;
        RECT 137.615 219.200 137.905 219.245 ;
        RECT 133.905 219.060 137.905 219.200 ;
        RECT 140.920 219.155 141.060 219.310 ;
        RECT 145.865 219.200 146.155 219.245 ;
        RECT 147.055 219.200 147.345 219.245 ;
        RECT 149.575 219.200 149.865 219.245 ;
        RECT 133.905 219.015 134.195 219.060 ;
        RECT 135.095 219.015 135.385 219.060 ;
        RECT 137.615 219.015 137.905 219.060 ;
        RECT 114.610 218.910 114.930 218.970 ;
        RECT 119.760 218.910 119.900 218.970 ;
        RECT 119.760 218.875 120.360 218.910 ;
        RECT 101.700 218.630 105.640 218.770 ;
        RECT 113.230 218.815 113.550 218.830 ;
        RECT 113.230 218.770 113.580 218.815 ;
        RECT 113.230 218.630 113.745 218.770 ;
        RECT 101.700 218.585 101.990 218.630 ;
        RECT 113.230 218.585 113.580 218.630 ;
        RECT 98.985 218.430 99.275 218.475 ;
        RECT 97.680 218.290 99.275 218.430 ;
        RECT 100.440 218.430 100.580 218.585 ;
        RECT 113.230 218.570 113.550 218.585 ;
        RECT 116.910 218.570 117.230 218.830 ;
        RECT 117.385 218.585 117.675 218.815 ;
        RECT 119.760 218.770 120.435 218.875 ;
        RECT 121.525 218.770 121.815 218.815 ;
        RECT 120.145 218.645 121.815 218.770 ;
        RECT 120.220 218.630 121.815 218.645 ;
        RECT 122.060 218.770 122.200 218.970 ;
        RECT 140.845 218.925 141.135 219.155 ;
        RECT 145.865 219.060 149.865 219.200 ;
        RECT 145.865 219.015 146.155 219.060 ;
        RECT 147.055 219.015 147.345 219.060 ;
        RECT 149.575 219.015 149.865 219.060 ;
        RECT 155.550 218.910 155.870 219.170 ;
        RECT 122.890 218.815 123.210 218.830 ;
        RECT 134.390 218.815 134.710 218.830 ;
        RECT 122.750 218.770 123.210 218.815 ;
        RECT 133.025 218.770 133.315 218.815 ;
        RECT 122.060 218.630 123.210 218.770 ;
        RECT 121.525 218.585 121.815 218.630 ;
        RECT 122.750 218.585 123.210 218.630 ;
        RECT 114.610 218.430 114.930 218.490 ;
        RECT 100.440 218.290 114.930 218.430 ;
        RECT 76.430 218.230 76.750 218.290 ;
        RECT 78.285 218.245 78.575 218.290 ;
        RECT 93.910 218.230 94.230 218.290 ;
        RECT 97.145 218.245 97.435 218.290 ;
        RECT 98.985 218.245 99.275 218.290 ;
        RECT 114.610 218.230 114.930 218.290 ;
        RECT 115.070 218.230 115.390 218.490 ;
        RECT 115.990 218.430 116.310 218.490 ;
        RECT 117.460 218.430 117.600 218.585 ;
        RECT 115.990 218.290 117.600 218.430 ;
        RECT 117.830 218.430 118.150 218.490 ;
        RECT 119.685 218.430 119.975 218.475 ;
        RECT 117.830 218.290 119.975 218.430 ;
        RECT 121.600 218.430 121.740 218.585 ;
        RECT 122.890 218.570 123.210 218.585 ;
        RECT 123.395 218.630 133.315 218.770 ;
        RECT 121.970 218.430 122.290 218.490 ;
        RECT 123.395 218.430 123.535 218.630 ;
        RECT 133.025 218.585 133.315 218.630 ;
        RECT 134.360 218.585 134.710 218.815 ;
        RECT 144.970 218.770 145.290 218.830 ;
        RECT 146.350 218.815 146.670 218.830 ;
        RECT 121.600 218.290 123.535 218.430 ;
        RECT 127.490 218.430 127.810 218.490 ;
        RECT 128.425 218.430 128.715 218.475 ;
        RECT 127.490 218.290 128.715 218.430 ;
        RECT 133.100 218.430 133.240 218.585 ;
        RECT 134.390 218.570 134.710 218.585 ;
        RECT 134.940 218.630 145.290 218.770 ;
        RECT 134.940 218.430 135.080 218.630 ;
        RECT 144.970 218.570 145.290 218.630 ;
        RECT 146.320 218.585 146.670 218.815 ;
        RECT 146.350 218.570 146.670 218.585 ;
        RECT 133.100 218.290 135.080 218.430 ;
        RECT 115.990 218.230 116.310 218.290 ;
        RECT 117.830 218.230 118.150 218.290 ;
        RECT 119.685 218.245 119.975 218.290 ;
        RECT 121.970 218.230 122.290 218.290 ;
        RECT 127.490 218.230 127.810 218.290 ;
        RECT 128.425 218.245 128.715 218.290 ;
        RECT 139.910 218.230 140.230 218.490 ;
        RECT 141.750 218.230 142.070 218.490 ;
        RECT 142.225 218.430 142.515 218.475 ;
        RECT 143.130 218.430 143.450 218.490 ;
        RECT 142.225 218.290 143.450 218.430 ;
        RECT 142.225 218.245 142.515 218.290 ;
        RECT 143.130 218.230 143.450 218.290 ;
        RECT 144.065 218.430 144.355 218.475 ;
        RECT 146.810 218.430 147.130 218.490 ;
        RECT 144.065 218.290 147.130 218.430 ;
        RECT 144.065 218.245 144.355 218.290 ;
        RECT 146.810 218.230 147.130 218.290 ;
        RECT 2.760 217.360 159.040 217.840 ;
        RECT 70.910 216.870 71.230 217.130 ;
        RECT 72.305 217.070 72.595 217.115 ;
        RECT 96.210 217.070 96.530 217.130 ;
        RECT 71.460 216.930 75.280 217.070 ;
        RECT 65.850 216.730 66.170 216.790 ;
        RECT 71.460 216.730 71.600 216.930 ;
        RECT 72.305 216.885 72.595 216.930 ;
        RECT 65.850 216.590 71.600 216.730 ;
        RECT 65.850 216.530 66.170 216.590 ;
        RECT 75.140 216.535 75.280 216.930 ;
        RECT 78.780 216.930 96.530 217.070 ;
        RECT 65.390 216.190 65.710 216.450 ;
        RECT 66.310 216.390 66.630 216.450 ;
        RECT 71.830 216.435 72.150 216.450 ;
        RECT 71.720 216.390 72.150 216.435 ;
        RECT 66.310 216.250 72.150 216.390 ;
        RECT 66.310 216.190 66.630 216.250 ;
        RECT 71.720 216.205 72.150 216.250 ;
        RECT 74.145 216.390 74.435 216.435 ;
        RECT 74.590 216.390 74.910 216.450 ;
        RECT 74.145 216.250 74.910 216.390 ;
        RECT 75.065 216.305 75.355 216.535 ;
        RECT 78.780 216.475 78.920 216.930 ;
        RECT 96.210 216.870 96.530 216.930 ;
        RECT 96.670 216.870 96.990 217.130 ;
        RECT 113.230 217.070 113.550 217.130 ;
        RECT 81.950 216.775 82.270 216.790 ;
        RECT 81.920 216.730 82.270 216.775 ;
        RECT 81.755 216.590 82.270 216.730 ;
        RECT 81.920 216.545 82.270 216.590 ;
        RECT 81.950 216.530 82.270 216.545 ;
        RECT 93.910 216.775 94.230 216.790 ;
        RECT 93.910 216.730 94.260 216.775 ;
        RECT 96.760 216.730 96.900 216.870 ;
        RECT 93.910 216.590 94.425 216.730 ;
        RECT 95.380 216.590 96.900 216.730 ;
        RECT 98.050 216.700 98.370 216.960 ;
        RECT 104.120 216.930 113.550 217.070 ;
        RECT 104.120 216.865 104.260 216.930 ;
        RECT 113.230 216.870 113.550 216.930 ;
        RECT 114.610 216.870 114.930 217.130 ;
        RECT 116.910 217.070 117.230 217.130 ;
        RECT 129.805 217.070 130.095 217.115 ;
        RECT 133.010 217.070 133.330 217.130 ;
        RECT 116.910 216.930 129.560 217.070 ;
        RECT 116.910 216.870 117.230 216.930 ;
        RECT 100.345 216.820 100.995 216.865 ;
        RECT 103.945 216.820 104.260 216.865 ;
        RECT 100.345 216.680 104.260 216.820 ;
        RECT 100.345 216.635 100.995 216.680 ;
        RECT 103.645 216.660 104.260 216.680 ;
        RECT 115.990 216.730 116.310 216.790 ;
        RECT 119.070 216.730 119.360 216.775 ;
        RECT 103.645 216.635 104.235 216.660 ;
        RECT 93.910 216.545 94.260 216.590 ;
        RECT 93.910 216.530 94.230 216.545 ;
        RECT 76.890 216.390 77.210 216.450 ;
        RECT 78.705 216.390 78.995 216.475 ;
        RECT 95.380 216.435 95.520 216.590 ;
        RECT 97.150 216.480 97.440 216.525 ;
        RECT 98.985 216.480 99.275 216.525 ;
        RECT 102.565 216.480 102.855 216.525 ;
        RECT 74.145 216.205 74.435 216.250 ;
        RECT 71.830 216.190 72.150 216.205 ;
        RECT 74.590 216.190 74.910 216.250 ;
        RECT 76.890 216.250 78.995 216.390 ;
        RECT 76.890 216.190 77.210 216.250 ;
        RECT 78.705 216.245 78.995 216.250 ;
        RECT 79.205 216.390 79.495 216.435 ;
        RECT 80.585 216.390 80.875 216.435 ;
        RECT 79.205 216.250 80.875 216.390 ;
        RECT 79.205 216.205 79.495 216.250 ;
        RECT 80.585 216.205 80.875 216.250 ;
        RECT 95.305 216.205 95.595 216.435 ;
        RECT 96.210 216.390 96.530 216.450 ;
        RECT 96.685 216.390 96.975 216.435 ;
        RECT 96.210 216.250 96.975 216.390 ;
        RECT 97.150 216.340 102.855 216.480 ;
        RECT 97.150 216.295 97.440 216.340 ;
        RECT 98.985 216.295 99.275 216.340 ;
        RECT 102.565 216.295 102.855 216.340 ;
        RECT 103.645 216.320 103.935 216.635 ;
        RECT 115.990 216.590 119.360 216.730 ;
        RECT 115.990 216.530 116.310 216.590 ;
        RECT 119.070 216.545 119.360 216.590 ;
        RECT 119.670 216.730 119.990 216.790 ;
        RECT 123.350 216.730 123.670 216.790 ;
        RECT 125.665 216.730 125.955 216.775 ;
        RECT 119.670 216.590 123.120 216.730 ;
        RECT 119.670 216.530 119.990 216.590 ;
        RECT 96.210 216.190 96.530 216.250 ;
        RECT 96.685 216.205 96.975 216.250 ;
        RECT 107.250 216.190 107.570 216.450 ;
        RECT 117.830 216.190 118.150 216.450 ;
        RECT 122.980 216.390 123.120 216.590 ;
        RECT 123.350 216.590 125.955 216.730 ;
        RECT 123.350 216.530 123.670 216.590 ;
        RECT 125.665 216.545 125.955 216.590 ;
        RECT 127.490 216.530 127.810 216.790 ;
        RECT 129.420 216.730 129.560 216.930 ;
        RECT 129.805 216.930 133.330 217.070 ;
        RECT 129.805 216.885 130.095 216.930 ;
        RECT 133.010 216.870 133.330 216.930 ;
        RECT 134.390 216.870 134.710 217.130 ;
        RECT 141.750 217.070 142.070 217.130 ;
        RECT 144.525 217.070 144.815 217.115 ;
        RECT 141.750 216.930 144.815 217.070 ;
        RECT 141.750 216.870 142.070 216.930 ;
        RECT 144.525 216.885 144.815 216.930 ;
        RECT 145.905 216.885 146.195 217.115 ;
        RECT 147.730 217.070 148.050 217.130 ;
        RECT 154.170 217.070 154.490 217.130 ;
        RECT 154.645 217.070 154.935 217.115 ;
        RECT 147.730 216.930 153.020 217.070 ;
        RECT 139.910 216.730 140.230 216.790 ;
        RECT 129.420 216.590 140.230 216.730 ;
        RECT 139.910 216.530 140.230 216.590 ;
        RECT 142.840 216.730 143.130 216.775 ;
        RECT 145.980 216.730 146.120 216.885 ;
        RECT 147.730 216.870 148.050 216.930 ;
        RECT 142.840 216.590 146.120 216.730 ;
        RECT 148.620 216.730 148.910 216.775 ;
        RECT 152.330 216.730 152.650 216.790 ;
        RECT 148.620 216.590 152.650 216.730 ;
        RECT 142.840 216.545 143.130 216.590 ;
        RECT 148.620 216.545 148.910 216.590 ;
        RECT 152.330 216.530 152.650 216.590 ;
        RECT 122.980 216.250 124.960 216.390 ;
        RECT 81.465 216.140 81.755 216.185 ;
        RECT 82.655 216.140 82.945 216.185 ;
        RECT 85.175 216.140 85.465 216.185 ;
        RECT 56.650 215.850 56.970 216.110 ;
        RECT 63.090 216.050 63.410 216.110 ;
        RECT 67.245 216.050 67.535 216.095 ;
        RECT 63.090 215.910 67.535 216.050 ;
        RECT 63.090 215.850 63.410 215.910 ;
        RECT 67.245 215.865 67.535 215.910 ;
        RECT 67.690 216.050 68.010 216.110 ;
        RECT 72.765 216.050 73.055 216.095 ;
        RECT 76.430 216.050 76.750 216.110 ;
        RECT 67.690 215.910 76.750 216.050 ;
        RECT 81.465 216.000 85.465 216.140 ;
        RECT 90.715 216.140 91.005 216.185 ;
        RECT 93.235 216.140 93.525 216.185 ;
        RECT 94.425 216.140 94.715 216.185 ;
        RECT 81.465 215.955 81.755 216.000 ;
        RECT 82.655 215.955 82.945 216.000 ;
        RECT 85.175 215.955 85.465 216.000 ;
        RECT 86.550 216.050 86.870 216.110 ;
        RECT 88.405 216.050 88.695 216.095 ;
        RECT 89.770 216.050 90.090 216.110 ;
        RECT 67.690 215.850 68.010 215.910 ;
        RECT 72.765 215.865 73.055 215.910 ;
        RECT 76.430 215.850 76.750 215.910 ;
        RECT 86.550 215.910 90.090 216.050 ;
        RECT 90.715 216.000 94.715 216.140 ;
        RECT 90.715 215.955 91.005 216.000 ;
        RECT 93.235 215.955 93.525 216.000 ;
        RECT 94.425 215.955 94.715 216.000 ;
        RECT 118.725 216.140 119.015 216.185 ;
        RECT 119.915 216.140 120.205 216.185 ;
        RECT 122.435 216.140 122.725 216.185 ;
        RECT 118.725 216.000 122.725 216.140 ;
        RECT 124.820 216.095 124.960 216.250 ;
        RECT 126.110 216.230 126.430 216.490 ;
        RECT 132.550 216.390 132.870 216.450 ;
        RECT 133.025 216.390 133.315 216.435 ;
        RECT 127.120 216.250 132.320 216.390 ;
        RECT 118.725 215.955 119.015 216.000 ;
        RECT 119.915 215.955 120.205 216.000 ;
        RECT 122.435 215.955 122.725 216.000 ;
        RECT 86.550 215.850 86.870 215.910 ;
        RECT 88.405 215.865 88.695 215.910 ;
        RECT 89.770 215.850 90.090 215.910 ;
        RECT 124.745 215.865 125.035 216.095 ;
        RECT 125.190 216.050 125.510 216.110 ;
        RECT 127.120 216.050 127.260 216.250 ;
        RECT 125.190 215.910 127.260 216.050 ;
        RECT 81.070 215.800 81.360 215.845 ;
        RECT 83.170 215.800 83.460 215.845 ;
        RECT 84.740 215.800 85.030 215.845 ;
        RECT 58.950 215.710 59.270 215.770 ;
        RECT 75.970 215.710 76.290 215.770 ;
        RECT 80.570 215.710 80.890 215.770 ;
        RECT 58.950 215.570 80.890 215.710 ;
        RECT 81.070 215.660 85.030 215.800 ;
        RECT 91.150 215.800 91.440 215.845 ;
        RECT 92.720 215.800 93.010 215.845 ;
        RECT 94.820 215.800 95.110 215.845 ;
        RECT 81.070 215.615 81.360 215.660 ;
        RECT 83.170 215.615 83.460 215.660 ;
        RECT 84.740 215.615 85.030 215.660 ;
        RECT 85.170 215.710 85.490 215.770 ;
        RECT 87.485 215.710 87.775 215.755 ;
        RECT 58.950 215.510 59.270 215.570 ;
        RECT 75.970 215.510 76.290 215.570 ;
        RECT 80.570 215.510 80.890 215.570 ;
        RECT 85.170 215.570 87.775 215.710 ;
        RECT 91.150 215.660 95.110 215.800 ;
        RECT 91.150 215.615 91.440 215.660 ;
        RECT 92.720 215.615 93.010 215.660 ;
        RECT 94.820 215.615 95.110 215.660 ;
        RECT 97.555 215.800 97.845 215.845 ;
        RECT 99.445 215.800 99.735 215.845 ;
        RECT 102.565 215.800 102.855 215.845 ;
        RECT 97.555 215.660 102.855 215.800 ;
        RECT 118.330 215.800 118.620 215.845 ;
        RECT 120.430 215.800 120.720 215.845 ;
        RECT 122.000 215.800 122.290 215.845 ;
        RECT 97.555 215.615 97.845 215.660 ;
        RECT 99.445 215.615 99.735 215.660 ;
        RECT 102.565 215.615 102.855 215.660 ;
        RECT 105.425 215.710 105.715 215.755 ;
        RECT 112.770 215.710 113.090 215.770 ;
        RECT 85.170 215.510 85.490 215.570 ;
        RECT 87.485 215.525 87.775 215.570 ;
        RECT 105.425 215.570 113.090 215.710 ;
        RECT 118.330 215.660 122.290 215.800 ;
        RECT 118.330 215.615 118.620 215.660 ;
        RECT 120.430 215.615 120.720 215.660 ;
        RECT 122.000 215.615 122.290 215.660 ;
        RECT 124.820 215.710 124.960 215.865 ;
        RECT 125.190 215.850 125.510 215.910 ;
        RECT 127.505 215.710 127.795 215.925 ;
        RECT 130.250 215.850 130.570 216.110 ;
        RECT 131.170 215.850 131.490 216.110 ;
        RECT 132.180 216.050 132.320 216.250 ;
        RECT 132.550 216.250 133.315 216.390 ;
        RECT 132.550 216.190 132.870 216.250 ;
        RECT 133.025 216.205 133.315 216.250 ;
        RECT 135.310 216.190 135.630 216.450 ;
        RECT 144.065 216.205 144.355 216.435 ;
        RECT 144.510 216.390 144.830 216.450 ;
        RECT 145.445 216.390 145.735 216.435 ;
        RECT 144.510 216.250 145.735 216.390 ;
        RECT 139.475 216.140 139.765 216.185 ;
        RECT 141.995 216.140 142.285 216.185 ;
        RECT 143.185 216.140 143.475 216.185 ;
        RECT 137.150 216.050 137.470 216.110 ;
        RECT 132.180 215.910 137.470 216.050 ;
        RECT 139.475 216.000 143.475 216.140 ;
        RECT 139.475 215.955 139.765 216.000 ;
        RECT 141.995 215.955 142.285 216.000 ;
        RECT 143.185 215.955 143.475 216.000 ;
        RECT 144.140 216.050 144.280 216.205 ;
        RECT 144.510 216.190 144.830 216.250 ;
        RECT 145.445 216.205 145.735 216.250 ;
        RECT 146.810 216.190 147.130 216.450 ;
        RECT 147.285 216.205 147.575 216.435 ;
        RECT 152.880 216.390 153.020 216.930 ;
        RECT 154.170 216.930 154.935 217.070 ;
        RECT 154.170 216.870 154.490 216.930 ;
        RECT 154.645 216.885 154.935 216.930 ;
        RECT 155.565 216.390 155.855 216.435 ;
        RECT 152.880 216.250 155.855 216.390 ;
        RECT 155.565 216.205 155.855 216.250 ;
        RECT 144.970 216.050 145.290 216.110 ;
        RECT 147.360 216.050 147.500 216.205 ;
        RECT 144.140 215.910 147.500 216.050 ;
        RECT 148.165 216.140 148.455 216.185 ;
        RECT 149.355 216.140 149.645 216.185 ;
        RECT 151.875 216.140 152.165 216.185 ;
        RECT 148.165 216.000 152.165 216.140 ;
        RECT 148.165 215.955 148.455 216.000 ;
        RECT 149.355 215.955 149.645 216.000 ;
        RECT 151.875 215.955 152.165 216.000 ;
        RECT 137.150 215.850 137.470 215.910 ;
        RECT 144.970 215.850 145.290 215.910 ;
        RECT 139.910 215.800 140.200 215.845 ;
        RECT 141.480 215.800 141.770 215.845 ;
        RECT 143.580 215.800 143.870 215.845 ;
        RECT 124.820 215.695 127.795 215.710 ;
        RECT 124.820 215.570 127.720 215.695 ;
        RECT 105.425 215.525 105.715 215.570 ;
        RECT 112.770 215.510 113.090 215.570 ;
        RECT 132.090 215.510 132.410 215.770 ;
        RECT 139.910 215.660 143.870 215.800 ;
        RECT 139.910 215.615 140.200 215.660 ;
        RECT 141.480 215.615 141.770 215.660 ;
        RECT 143.580 215.615 143.870 215.660 ;
        RECT 147.770 215.800 148.060 215.845 ;
        RECT 149.870 215.800 150.160 215.845 ;
        RECT 151.440 215.800 151.730 215.845 ;
        RECT 147.770 215.660 151.730 215.800 ;
        RECT 147.770 215.615 148.060 215.660 ;
        RECT 149.870 215.615 150.160 215.660 ;
        RECT 151.440 215.615 151.730 215.660 ;
        RECT 154.185 215.710 154.475 215.755 ;
        RECT 155.550 215.710 155.870 215.770 ;
        RECT 154.185 215.570 155.870 215.710 ;
        RECT 154.185 215.525 154.475 215.570 ;
        RECT 155.550 215.510 155.870 215.570 ;
        RECT 1.000 214.640 158.240 215.120 ;
        RECT 55.730 214.150 56.050 214.410 ;
        RECT 58.505 214.350 58.795 214.395 ;
        RECT 62.170 214.350 62.490 214.410 ;
        RECT 58.505 214.210 62.490 214.350 ;
        RECT 58.505 214.165 58.795 214.210 ;
        RECT 62.170 214.150 62.490 214.210 ;
        RECT 65.390 214.350 65.710 214.410 ;
        RECT 84.265 214.350 84.555 214.395 ;
        RECT 107.250 214.350 107.570 214.410 ;
        RECT 65.390 214.210 107.570 214.350 ;
        RECT 65.390 214.150 65.710 214.210 ;
        RECT 84.265 214.165 84.555 214.210 ;
        RECT 107.250 214.150 107.570 214.210 ;
        RECT 109.090 214.350 109.410 214.410 ;
        RECT 116.925 214.350 117.215 214.395 ;
        RECT 132.090 214.350 132.410 214.410 ;
        RECT 109.090 214.210 117.215 214.350 ;
        RECT 109.090 214.150 109.410 214.210 ;
        RECT 116.925 214.165 117.215 214.210 ;
        RECT 127.580 214.210 132.410 214.350 ;
        RECT 122.470 214.100 122.760 214.145 ;
        RECT 124.570 214.100 124.860 214.145 ;
        RECT 126.140 214.100 126.430 214.145 ;
        RECT 63.090 214.010 63.410 214.070 ;
        RECT 63.565 214.010 63.855 214.055 ;
        RECT 63.090 213.870 63.855 214.010 ;
        RECT 63.090 213.810 63.410 213.870 ;
        RECT 63.565 213.825 63.855 213.870 ;
        RECT 66.770 214.010 67.090 214.070 ;
        RECT 76.890 214.010 77.210 214.070 ;
        RECT 120.145 214.010 120.435 214.055 ;
        RECT 120.590 214.010 120.910 214.070 ;
        RECT 66.770 213.870 73.900 214.010 ;
        RECT 66.770 213.810 67.090 213.870 ;
        RECT 59.885 213.670 60.175 213.715 ;
        RECT 56.280 213.530 60.175 213.670 ;
        RECT 56.280 213.375 56.420 213.530 ;
        RECT 59.885 213.485 60.175 213.530 ;
        RECT 61.265 213.670 61.555 213.715 ;
        RECT 66.860 213.670 67.000 213.810 ;
        RECT 73.760 213.715 73.900 213.870 ;
        RECT 61.265 213.530 67.000 213.670 ;
        RECT 73.685 213.670 73.975 213.715 ;
        RECT 74.590 213.670 74.910 213.730 ;
        RECT 73.685 213.530 74.910 213.670 ;
        RECT 61.265 213.485 61.555 213.530 ;
        RECT 73.685 213.485 73.975 213.530 ;
        RECT 74.590 213.470 74.910 213.530 ;
        RECT 75.050 213.670 75.370 213.730 ;
        RECT 75.985 213.670 76.275 213.885 ;
        RECT 76.890 213.870 79.420 214.010 ;
        RECT 76.890 213.810 77.210 213.870 ;
        RECT 75.050 213.655 76.275 213.670 ;
        RECT 75.050 213.530 76.200 213.655 ;
        RECT 75.050 213.470 75.370 213.530 ;
        RECT 67.230 213.405 67.550 213.465 ;
        RECT 79.280 213.450 79.420 213.870 ;
        RECT 97.680 213.870 119.440 214.010 ;
        RECT 84.710 213.670 85.030 213.730 ;
        RECT 84.710 213.530 92.300 213.670 ;
        RECT 84.710 213.470 85.030 213.530 ;
        RECT 68.395 213.405 68.685 213.450 ;
        RECT 56.205 213.145 56.495 213.375 ;
        RECT 58.965 213.330 59.255 213.375 ;
        RECT 62.630 213.330 62.950 213.390 ;
        RECT 58.965 213.190 62.950 213.330 ;
        RECT 58.965 213.145 59.255 213.190 ;
        RECT 62.630 213.130 62.950 213.190 ;
        RECT 60.790 212.790 61.110 213.050 ;
        RECT 61.710 212.990 62.030 213.050 ;
        RECT 63.565 212.990 63.855 213.205 ;
        RECT 64.930 213.130 65.250 213.390 ;
        RECT 65.390 213.330 65.710 213.390 ;
        RECT 66.785 213.330 67.075 213.375 ;
        RECT 65.390 213.190 67.075 213.330 ;
        RECT 67.230 213.265 68.685 213.405 ;
        RECT 67.230 213.205 67.550 213.265 ;
        RECT 68.395 213.220 68.685 213.265 ;
        RECT 71.385 213.330 71.675 213.450 ;
        RECT 75.970 213.330 76.290 213.390 ;
        RECT 71.385 213.220 76.290 213.330 ;
        RECT 71.460 213.190 76.290 213.220 ;
        RECT 65.390 213.130 65.710 213.190 ;
        RECT 66.785 213.145 67.075 213.190 ;
        RECT 75.970 213.130 76.290 213.190 ;
        RECT 76.430 213.330 76.750 213.390 ;
        RECT 77.825 213.330 78.115 213.375 ;
        RECT 78.270 213.330 78.590 213.390 ;
        RECT 76.430 213.190 77.580 213.330 ;
        RECT 76.430 213.130 76.750 213.190 ;
        RECT 67.690 212.990 68.010 213.050 ;
        RECT 61.710 212.850 68.010 212.990 ;
        RECT 61.710 212.790 62.030 212.850 ;
        RECT 67.690 212.790 68.010 212.850 ;
        RECT 70.910 212.790 71.230 213.050 ;
        RECT 74.605 212.990 74.895 213.035 ;
        RECT 76.890 212.990 77.210 213.050 ;
        RECT 74.605 212.850 77.210 212.990 ;
        RECT 77.440 212.990 77.580 213.190 ;
        RECT 77.825 213.190 78.590 213.330 ;
        RECT 79.205 213.220 79.495 213.450 ;
        RECT 81.490 213.205 81.810 213.465 ;
        RECT 92.160 213.375 92.300 213.530 ;
        RECT 90.705 213.330 90.995 213.375 ;
        RECT 77.825 213.145 78.115 213.190 ;
        RECT 78.270 213.130 78.590 213.190 ;
        RECT 90.705 213.190 91.840 213.330 ;
        RECT 90.705 213.145 90.995 213.190 ;
        RECT 86.550 212.990 86.870 213.050 ;
        RECT 77.440 212.850 86.870 212.990 ;
        RECT 74.605 212.805 74.895 212.850 ;
        RECT 76.890 212.790 77.210 212.850 ;
        RECT 86.550 212.790 86.870 212.850 ;
        RECT 91.150 212.790 91.470 213.050 ;
        RECT 91.700 212.990 91.840 213.190 ;
        RECT 92.085 213.145 92.375 213.375 ;
        RECT 97.680 212.990 97.820 213.870 ;
        RECT 98.050 213.670 98.370 213.730 ;
        RECT 104.490 213.670 104.810 213.730 ;
        RECT 98.050 213.530 104.810 213.670 ;
        RECT 98.050 213.470 98.370 213.530 ;
        RECT 104.490 213.470 104.810 213.530 ;
        RECT 104.965 213.485 105.255 213.715 ;
        RECT 105.410 213.670 105.730 213.730 ;
        RECT 106.345 213.670 106.635 213.715 ;
        RECT 105.410 213.530 106.635 213.670 ;
        RECT 105.040 213.330 105.180 213.485 ;
        RECT 105.410 213.470 105.730 213.530 ;
        RECT 106.345 213.485 106.635 213.530 ;
        RECT 109.090 213.470 109.410 213.730 ;
        RECT 112.770 213.470 113.090 213.730 ;
        RECT 115.545 213.670 115.835 213.715 ;
        RECT 117.370 213.670 117.690 213.730 ;
        RECT 119.300 213.670 119.440 213.870 ;
        RECT 120.145 213.870 120.910 214.010 ;
        RECT 122.470 213.960 126.430 214.100 ;
        RECT 122.470 213.915 122.760 213.960 ;
        RECT 124.570 213.915 124.860 213.960 ;
        RECT 126.140 213.915 126.430 213.960 ;
        RECT 120.145 213.825 120.435 213.870 ;
        RECT 120.590 213.810 120.910 213.870 ;
        RECT 122.865 213.760 123.155 213.805 ;
        RECT 124.055 213.760 124.345 213.805 ;
        RECT 126.575 213.760 126.865 213.805 ;
        RECT 115.545 213.530 117.690 213.670 ;
        RECT 115.545 213.485 115.835 213.530 ;
        RECT 117.370 213.470 117.690 213.530 ;
        RECT 117.920 213.530 118.980 213.670 ;
        RECT 119.300 213.530 121.280 213.670 ;
        RECT 111.850 213.330 112.170 213.390 ;
        RECT 105.040 213.190 115.760 213.330 ;
        RECT 111.850 213.130 112.170 213.190 ;
        RECT 91.700 212.850 97.820 212.990 ;
        RECT 99.430 212.990 99.750 213.050 ;
        RECT 102.205 212.990 102.495 213.035 ;
        RECT 99.430 212.850 102.495 212.990 ;
        RECT 99.430 212.790 99.750 212.850 ;
        RECT 102.205 212.805 102.495 212.850 ;
        RECT 104.030 212.790 104.350 213.050 ;
        RECT 104.505 212.990 104.795 213.035 ;
        RECT 105.870 212.990 106.190 213.050 ;
        RECT 104.505 212.850 106.190 212.990 ;
        RECT 104.505 212.805 104.795 212.850 ;
        RECT 105.870 212.790 106.190 212.850 ;
        RECT 107.250 212.990 107.570 213.050 ;
        RECT 110.025 212.990 110.315 213.035 ;
        RECT 107.250 212.850 110.315 212.990 ;
        RECT 107.250 212.790 107.570 212.850 ;
        RECT 110.025 212.805 110.315 212.850 ;
        RECT 113.690 212.990 114.010 213.050 ;
        RECT 115.070 212.990 115.390 213.050 ;
        RECT 113.690 212.850 115.390 212.990 ;
        RECT 115.620 212.990 115.760 213.190 ;
        RECT 115.990 213.130 116.310 213.390 ;
        RECT 117.920 213.330 118.060 213.530 ;
        RECT 116.540 213.190 118.060 213.330 ;
        RECT 116.540 212.990 116.680 213.190 ;
        RECT 118.305 213.145 118.595 213.375 ;
        RECT 118.840 213.330 118.980 213.530 ;
        RECT 119.670 213.330 119.990 213.390 ;
        RECT 118.840 213.190 119.990 213.330 ;
        RECT 115.620 212.850 116.680 212.990 ;
        RECT 113.690 212.790 114.010 212.850 ;
        RECT 115.070 212.790 115.390 212.850 ;
        RECT 117.370 212.790 117.690 213.050 ;
        RECT 118.380 212.990 118.520 213.145 ;
        RECT 119.670 213.130 119.990 213.190 ;
        RECT 119.225 212.990 119.515 213.035 ;
        RECT 118.380 212.850 119.515 212.990 ;
        RECT 121.140 212.990 121.280 213.530 ;
        RECT 121.970 213.470 122.290 213.730 ;
        RECT 122.865 213.620 126.865 213.760 ;
        RECT 122.865 213.575 123.155 213.620 ;
        RECT 124.055 213.575 124.345 213.620 ;
        RECT 126.575 213.575 126.865 213.620 ;
        RECT 121.525 213.330 121.815 213.375 ;
        RECT 122.430 213.330 122.750 213.390 ;
        RECT 121.525 213.190 122.750 213.330 ;
        RECT 121.525 213.145 121.815 213.190 ;
        RECT 122.430 213.130 122.750 213.190 ;
        RECT 123.320 213.330 123.610 213.375 ;
        RECT 127.580 213.330 127.720 214.210 ;
        RECT 132.090 214.150 132.410 214.210 ;
        RECT 143.130 214.150 143.450 214.410 ;
        RECT 145.890 214.150 146.210 214.410 ;
        RECT 146.350 214.150 146.670 214.410 ;
        RECT 152.330 214.150 152.650 214.410 ;
        RECT 154.630 214.010 154.950 214.070 ;
        RECT 123.320 213.190 127.720 213.330 ;
        RECT 128.500 213.870 154.950 214.010 ;
        RECT 123.320 213.145 123.610 213.190 ;
        RECT 128.500 212.990 128.640 213.870 ;
        RECT 154.630 213.810 154.950 213.870 ;
        RECT 132.105 213.670 132.395 213.715 ;
        RECT 128.960 213.530 132.395 213.670 ;
        RECT 128.960 213.035 129.100 213.530 ;
        RECT 132.105 213.485 132.395 213.530 ;
        RECT 137.150 213.670 137.470 213.730 ;
        RECT 139.925 213.670 140.215 213.715 ;
        RECT 137.150 213.530 140.215 213.670 ;
        RECT 137.150 213.470 137.470 213.530 ;
        RECT 139.925 213.485 140.215 213.530 ;
        RECT 130.250 213.330 130.570 213.390 ;
        RECT 133.025 213.330 133.315 213.375 ;
        RECT 130.250 213.190 133.315 213.330 ;
        RECT 130.250 213.130 130.570 213.190 ;
        RECT 133.025 213.145 133.315 213.190 ;
        RECT 133.930 213.130 134.250 213.390 ;
        RECT 144.050 213.330 144.370 213.390 ;
        RECT 144.985 213.330 145.275 213.375 ;
        RECT 144.050 213.190 145.275 213.330 ;
        RECT 144.050 213.130 144.370 213.190 ;
        RECT 144.985 213.145 145.275 213.190 ;
        RECT 147.270 213.130 147.590 213.390 ;
        RECT 152.790 213.330 153.110 213.390 ;
        RECT 153.265 213.330 153.555 213.375 ;
        RECT 152.790 213.190 153.555 213.330 ;
        RECT 152.790 213.130 153.110 213.190 ;
        RECT 153.265 213.145 153.555 213.190 ;
        RECT 121.140 212.850 128.640 212.990 ;
        RECT 119.225 212.805 119.515 212.850 ;
        RECT 128.885 212.805 129.175 213.035 ;
        RECT 129.330 212.790 129.650 213.050 ;
        RECT 2.760 211.920 159.040 212.400 ;
        RECT 57.570 211.630 57.890 211.690 ;
        RECT 60.345 211.630 60.635 211.675 ;
        RECT 57.570 211.490 60.635 211.630 ;
        RECT 57.570 211.430 57.890 211.490 ;
        RECT 60.345 211.445 60.635 211.490 ;
        RECT 61.710 211.430 62.030 211.690 ;
        RECT 64.470 211.630 64.790 211.690 ;
        RECT 65.865 211.630 66.155 211.675 ;
        RECT 67.230 211.630 67.550 211.690 ;
        RECT 64.470 211.490 67.550 211.630 ;
        RECT 64.470 211.430 64.790 211.490 ;
        RECT 65.865 211.445 66.155 211.490 ;
        RECT 67.230 211.430 67.550 211.490 ;
        RECT 67.690 211.430 68.010 211.690 ;
        RECT 69.070 211.630 69.390 211.690 ;
        RECT 71.370 211.630 71.690 211.690 ;
        RECT 69.070 211.490 71.690 211.630 ;
        RECT 69.070 211.430 69.390 211.490 ;
        RECT 71.370 211.430 71.690 211.490 ;
        RECT 72.290 211.630 72.610 211.690 ;
        RECT 81.950 211.630 82.270 211.690 ;
        RECT 110.485 211.630 110.775 211.675 ;
        RECT 72.290 211.490 81.720 211.630 ;
        RECT 72.290 211.430 72.610 211.490 ;
        RECT 11.570 211.290 11.890 211.350 ;
        RECT 14.850 211.290 15.140 211.335 ;
        RECT 19.390 211.290 19.710 211.350 ;
        RECT 56.650 211.290 56.970 211.350 ;
        RECT 11.570 211.150 15.140 211.290 ;
        RECT 11.570 211.090 11.890 211.150 ;
        RECT 14.850 211.105 15.140 211.150 ;
        RECT 16.260 211.150 56.970 211.290 ;
        RECT 16.260 210.995 16.400 211.150 ;
        RECT 19.390 211.090 19.710 211.150 ;
        RECT 56.650 211.090 56.970 211.150 ;
        RECT 58.965 211.290 59.255 211.335 ;
        RECT 60.790 211.290 61.110 211.350 ;
        RECT 61.265 211.290 61.555 211.335 ;
        RECT 64.025 211.290 64.315 211.335 ;
        RECT 58.965 211.150 63.655 211.290 ;
        RECT 58.965 211.105 59.255 211.150 ;
        RECT 60.790 211.090 61.110 211.150 ;
        RECT 61.265 211.105 61.555 211.150 ;
        RECT 16.185 210.765 16.475 210.995 ;
        RECT 17.090 210.750 17.410 211.010 ;
        RECT 63.515 210.990 63.655 211.150 ;
        RECT 64.025 211.150 67.000 211.290 ;
        RECT 64.025 211.105 64.315 211.150 ;
        RECT 66.860 211.010 67.000 211.150 ;
        RECT 63.515 210.950 63.780 210.990 ;
        RECT 64.945 210.950 65.235 210.995 ;
        RECT 63.515 210.850 65.235 210.950 ;
        RECT 63.640 210.810 65.235 210.850 ;
        RECT 64.945 210.765 65.235 210.810 ;
        RECT 66.770 210.950 67.090 211.010 ;
        RECT 67.780 210.995 67.920 211.430 ;
        RECT 69.990 211.290 70.310 211.350 ;
        RECT 69.990 211.150 74.820 211.290 ;
        RECT 69.990 211.090 70.310 211.150 ;
        RECT 67.340 210.950 67.630 210.995 ;
        RECT 66.770 210.810 67.630 210.950 ;
        RECT 67.780 210.810 68.120 210.995 ;
        RECT 11.595 210.700 11.885 210.745 ;
        RECT 14.115 210.700 14.405 210.745 ;
        RECT 15.305 210.700 15.595 210.745 ;
        RECT 11.595 210.560 15.595 210.700 ;
        RECT 11.595 210.515 11.885 210.560 ;
        RECT 14.115 210.515 14.405 210.560 ;
        RECT 15.305 210.515 15.595 210.560 ;
        RECT 57.125 210.610 57.415 210.655 ;
        RECT 63.090 210.610 63.410 210.670 ;
        RECT 57.125 210.470 63.410 210.610 ;
        RECT 65.020 210.610 65.160 210.765 ;
        RECT 66.770 210.750 67.090 210.810 ;
        RECT 67.340 210.765 67.630 210.810 ;
        RECT 67.830 210.765 68.120 210.810 ;
        RECT 70.465 210.950 70.755 210.995 ;
        RECT 70.910 210.950 71.230 211.010 ;
        RECT 70.465 210.810 71.230 210.950 ;
        RECT 70.465 210.765 70.755 210.810 ;
        RECT 70.910 210.750 71.230 210.810 ;
        RECT 71.830 210.750 72.150 211.010 ;
        RECT 72.765 210.935 73.055 211.150 ;
        RECT 74.680 211.055 74.820 211.150 ;
        RECT 75.985 211.055 76.275 211.100 ;
        RECT 74.680 210.915 76.275 211.055 ;
        RECT 75.510 210.750 75.830 210.915 ;
        RECT 75.985 210.870 76.275 210.915 ;
        RECT 76.890 211.055 77.210 211.115 ;
        RECT 78.270 211.055 78.590 211.115 ;
        RECT 76.890 210.915 78.590 211.055 ;
        RECT 81.580 210.995 81.720 211.490 ;
        RECT 81.950 211.490 100.120 211.630 ;
        RECT 81.950 211.430 82.270 211.490 ;
        RECT 99.980 211.460 100.120 211.490 ;
        RECT 100.900 211.490 110.775 211.630 ;
        RECT 100.900 211.460 101.040 211.490 ;
        RECT 87.010 211.290 87.330 211.350 ;
        RECT 98.970 211.290 99.290 211.350 ;
        RECT 99.980 211.320 101.040 211.460 ;
        RECT 110.485 211.445 110.775 211.490 ;
        RECT 113.690 211.430 114.010 211.690 ;
        RECT 116.450 211.630 116.770 211.690 ;
        RECT 116.925 211.630 117.215 211.675 ;
        RECT 116.450 211.490 117.215 211.630 ;
        RECT 116.450 211.430 116.770 211.490 ;
        RECT 116.925 211.445 117.215 211.490 ;
        RECT 121.510 211.630 121.830 211.690 ;
        RECT 127.030 211.630 127.350 211.690 ;
        RECT 129.330 211.630 129.650 211.690 ;
        RECT 121.510 211.490 129.650 211.630 ;
        RECT 121.510 211.430 121.830 211.490 ;
        RECT 87.010 211.150 99.290 211.290 ;
        RECT 84.710 211.030 85.030 211.090 ;
        RECT 85.180 211.030 85.470 211.075 ;
        RECT 76.890 210.855 77.210 210.915 ;
        RECT 78.270 210.855 78.590 210.915 ;
        RECT 81.505 210.765 81.795 210.995 ;
        RECT 84.710 210.890 85.470 211.030 ;
        RECT 84.710 210.830 85.030 210.890 ;
        RECT 85.180 210.845 85.470 210.890 ;
        RECT 85.630 210.950 85.950 211.010 ;
        RECT 86.105 210.950 86.395 210.995 ;
        RECT 85.630 210.810 86.395 210.950 ;
        RECT 86.550 210.870 86.870 211.130 ;
        RECT 87.010 211.090 87.330 211.150 ;
        RECT 98.970 211.090 99.290 211.150 ;
        RECT 100.365 211.120 100.655 211.165 ;
        RECT 98.065 210.950 98.355 210.995 ;
        RECT 85.630 210.750 85.950 210.810 ;
        RECT 86.105 210.765 86.395 210.810 ;
        RECT 88.940 210.810 98.355 210.950 ;
        RECT 71.920 210.610 72.060 210.750 ;
        RECT 57.125 210.425 57.415 210.470 ;
        RECT 63.090 210.410 63.410 210.470 ;
        RECT 63.550 210.440 63.870 210.500 ;
        RECT 64.025 210.440 64.315 210.485 ;
        RECT 65.020 210.470 72.060 210.610 ;
        RECT 73.685 210.610 73.975 210.655 ;
        RECT 77.350 210.610 77.670 210.670 ;
        RECT 73.685 210.470 77.670 210.610 ;
        RECT 12.030 210.360 12.320 210.405 ;
        RECT 13.600 210.360 13.890 210.405 ;
        RECT 15.700 210.360 15.990 210.405 ;
        RECT 9.270 210.070 9.590 210.330 ;
        RECT 12.030 210.220 15.990 210.360 ;
        RECT 12.030 210.175 12.320 210.220 ;
        RECT 13.600 210.175 13.890 210.220 ;
        RECT 15.700 210.175 15.990 210.220 ;
        RECT 20.325 210.270 20.615 210.315 ;
        RECT 20.770 210.270 21.090 210.330 ;
        RECT 20.325 210.130 21.090 210.270 ;
        RECT 20.325 210.085 20.615 210.130 ;
        RECT 20.770 210.070 21.090 210.130 ;
        RECT 58.950 209.820 59.270 210.080 ;
        RECT 59.870 210.070 60.190 210.330 ;
        RECT 63.550 210.300 64.315 210.440 ;
        RECT 69.160 210.330 69.300 210.470 ;
        RECT 73.685 210.425 73.975 210.470 ;
        RECT 77.350 210.410 77.670 210.470 ;
        RECT 77.810 210.610 78.130 210.670 ;
        RECT 78.285 210.610 78.575 210.655 ;
        RECT 82.425 210.610 82.715 210.655 ;
        RECT 82.870 210.610 83.190 210.670 ;
        RECT 77.810 210.470 82.180 210.610 ;
        RECT 77.810 210.410 78.130 210.470 ;
        RECT 78.285 210.425 78.575 210.470 ;
        RECT 63.550 210.240 63.870 210.300 ;
        RECT 64.025 210.270 64.315 210.300 ;
        RECT 64.930 210.270 65.250 210.330 ;
        RECT 64.025 210.255 65.250 210.270 ;
        RECT 64.100 210.130 65.250 210.255 ;
        RECT 64.930 210.070 65.250 210.130 ;
        RECT 69.070 210.070 69.390 210.330 ;
        RECT 74.130 210.270 74.450 210.330 ;
        RECT 80.585 210.270 80.875 210.315 ;
        RECT 74.130 210.130 80.875 210.270 ;
        RECT 82.040 210.270 82.180 210.470 ;
        RECT 82.425 210.470 83.190 210.610 ;
        RECT 82.425 210.425 82.715 210.470 ;
        RECT 82.870 210.410 83.190 210.470 ;
        RECT 84.250 210.410 84.570 210.670 ;
        RECT 88.940 210.610 89.080 210.810 ;
        RECT 98.065 210.765 98.355 210.810 ;
        RECT 99.430 210.950 99.750 211.010 ;
        RECT 99.980 210.980 100.655 211.120 ;
        RECT 101.270 211.090 101.590 211.350 ;
        RECT 101.730 211.290 102.050 211.350 ;
        RECT 101.730 211.150 103.800 211.290 ;
        RECT 101.730 211.090 102.050 211.150 ;
        RECT 103.660 210.995 103.800 211.150 ;
        RECT 99.980 210.950 100.120 210.980 ;
        RECT 99.430 210.810 100.120 210.950 ;
        RECT 100.365 210.935 100.655 210.980 ;
        RECT 102.205 210.950 102.495 210.995 ;
        RECT 103.125 210.950 103.415 210.995 ;
        RECT 102.205 210.810 103.415 210.950 ;
        RECT 99.430 210.750 99.750 210.810 ;
        RECT 102.205 210.765 102.495 210.810 ;
        RECT 103.125 210.765 103.415 210.810 ;
        RECT 103.585 210.765 103.875 210.995 ;
        RECT 107.250 210.920 107.570 211.180 ;
        RECT 108.170 211.090 108.490 211.350 ;
        RECT 108.695 211.120 108.985 211.165 ;
        RECT 109.550 211.120 109.870 211.180 ;
        RECT 108.185 210.935 108.475 211.090 ;
        RECT 108.695 210.980 109.870 211.120 ;
        RECT 111.390 211.090 111.710 211.350 ;
        RECT 122.890 211.290 123.210 211.350 ;
        RECT 115.620 211.150 123.210 211.290 ;
        RECT 108.695 210.935 108.985 210.980 ;
        RECT 109.550 210.920 109.870 210.980 ;
        RECT 111.850 210.830 112.170 211.090 ;
        RECT 112.310 211.030 112.630 211.090 ;
        RECT 112.785 211.030 113.075 211.075 ;
        RECT 112.310 210.890 113.075 211.030 ;
        RECT 115.620 210.995 115.760 211.150 ;
        RECT 122.890 211.090 123.210 211.150 ;
        RECT 123.725 211.120 124.015 211.165 ;
        RECT 124.360 211.120 124.500 211.490 ;
        RECT 127.030 211.430 127.350 211.490 ;
        RECT 129.330 211.430 129.650 211.490 ;
        RECT 112.310 210.830 112.630 210.890 ;
        RECT 112.785 210.845 113.075 210.890 ;
        RECT 115.545 210.765 115.835 210.995 ;
        RECT 85.720 210.470 89.080 210.610 ;
        RECT 90.230 210.610 90.550 210.670 ;
        RECT 96.210 210.610 96.530 210.670 ;
        RECT 97.130 210.610 97.450 210.670 ;
        RECT 90.230 210.470 97.450 210.610 ;
        RECT 85.720 210.270 85.860 210.470 ;
        RECT 90.230 210.410 90.550 210.470 ;
        RECT 96.210 210.410 96.530 210.470 ;
        RECT 97.130 210.410 97.450 210.470 ;
        RECT 98.985 210.610 99.275 210.655 ;
        RECT 103.200 210.610 103.340 210.765 ;
        RECT 115.990 210.750 116.310 211.010 ;
        RECT 121.050 210.950 121.370 211.010 ;
        RECT 122.445 210.950 122.735 210.995 ;
        RECT 121.050 210.810 122.735 210.950 ;
        RECT 123.725 210.980 124.500 211.120 ;
        RECT 123.725 210.935 124.015 210.980 ;
        RECT 121.050 210.750 121.370 210.810 ;
        RECT 122.445 210.765 122.735 210.810 ;
        RECT 134.865 210.765 135.155 210.995 ;
        RECT 123.325 210.700 123.615 210.745 ;
        RECT 124.515 210.700 124.805 210.745 ;
        RECT 127.035 210.700 127.325 210.745 ;
        RECT 104.030 210.610 104.350 210.670 ;
        RECT 105.410 210.610 105.730 210.670 ;
        RECT 98.985 210.470 102.880 210.610 ;
        RECT 103.200 210.470 105.730 210.610 ;
        RECT 98.985 210.425 99.275 210.470 ;
        RECT 82.040 210.130 85.860 210.270 ;
        RECT 99.445 210.270 99.735 210.315 ;
        RECT 100.350 210.270 100.670 210.330 ;
        RECT 99.445 210.130 100.670 210.270 ;
        RECT 102.740 210.270 102.880 210.470 ;
        RECT 104.030 210.410 104.350 210.470 ;
        RECT 105.410 210.410 105.730 210.470 ;
        RECT 106.345 210.610 106.635 210.655 ;
        RECT 109.090 210.610 109.410 210.670 ;
        RECT 113.230 210.610 113.550 210.670 ;
        RECT 106.345 210.470 109.410 210.610 ;
        RECT 106.345 210.425 106.635 210.470 ;
        RECT 109.090 210.410 109.410 210.470 ;
        RECT 111.940 210.470 113.550 210.610 ;
        RECT 123.325 210.560 127.325 210.700 ;
        RECT 123.325 210.515 123.615 210.560 ;
        RECT 124.515 210.515 124.805 210.560 ;
        RECT 127.035 210.515 127.325 210.560 ;
        RECT 129.345 210.610 129.635 210.655 ;
        RECT 134.940 210.610 135.080 210.765 ;
        RECT 103.570 210.270 103.890 210.330 ;
        RECT 102.740 210.130 103.890 210.270 ;
        RECT 71.370 209.820 71.690 210.080 ;
        RECT 74.130 210.070 74.450 210.130 ;
        RECT 80.585 210.085 80.875 210.130 ;
        RECT 99.445 210.085 99.735 210.130 ;
        RECT 100.350 210.070 100.670 210.130 ;
        RECT 103.570 210.070 103.890 210.130 ;
        RECT 104.490 210.070 104.810 210.330 ;
        RECT 106.790 210.270 107.110 210.330 ;
        RECT 109.565 210.270 109.855 210.315 ;
        RECT 106.790 210.130 109.855 210.270 ;
        RECT 106.790 210.070 107.110 210.130 ;
        RECT 109.565 210.085 109.855 210.130 ;
        RECT 110.655 210.020 110.945 210.065 ;
        RECT 111.940 210.020 112.080 210.470 ;
        RECT 113.230 210.410 113.550 210.470 ;
        RECT 129.345 210.470 135.080 210.610 ;
        RECT 129.345 210.425 129.635 210.470 ;
        RECT 122.930 210.360 123.220 210.405 ;
        RECT 125.030 210.360 125.320 210.405 ;
        RECT 126.600 210.360 126.890 210.405 ;
        RECT 112.310 210.270 112.630 210.330 ;
        RECT 112.785 210.270 113.075 210.315 ;
        RECT 112.310 210.130 113.075 210.270 ;
        RECT 122.930 210.220 126.890 210.360 ;
        RECT 122.930 210.175 123.220 210.220 ;
        RECT 125.030 210.175 125.320 210.220 ;
        RECT 126.600 210.175 126.890 210.220 ;
        RECT 128.410 210.270 128.730 210.330 ;
        RECT 132.105 210.270 132.395 210.315 ;
        RECT 112.310 210.070 112.630 210.130 ;
        RECT 112.785 210.085 113.075 210.130 ;
        RECT 128.410 210.130 132.395 210.270 ;
        RECT 128.410 210.070 128.730 210.130 ;
        RECT 132.105 210.085 132.395 210.130 ;
        RECT 110.655 209.880 112.080 210.020 ;
        RECT 110.655 209.835 110.945 209.880 ;
        RECT 1.000 209.200 158.240 209.680 ;
        RECT 61.710 208.910 62.030 208.970 ;
        RECT 70.925 208.910 71.215 208.955 ;
        RECT 72.750 208.910 73.070 208.970 ;
        RECT 81.490 208.910 81.810 208.970 ;
        RECT 84.710 208.910 85.030 208.970 ;
        RECT 61.710 208.770 73.070 208.910 ;
        RECT 61.710 208.710 62.030 208.770 ;
        RECT 70.925 208.725 71.215 208.770 ;
        RECT 72.750 208.710 73.070 208.770 ;
        RECT 74.680 208.770 81.810 208.910 ;
        RECT 19.890 208.660 20.180 208.705 ;
        RECT 21.990 208.660 22.280 208.705 ;
        RECT 23.560 208.660 23.850 208.705 ;
        RECT 19.890 208.520 23.850 208.660 ;
        RECT 19.890 208.475 20.180 208.520 ;
        RECT 21.990 208.475 22.280 208.520 ;
        RECT 23.560 208.475 23.850 208.520 ;
        RECT 33.205 208.570 33.495 208.615 ;
        RECT 74.680 208.570 74.820 208.770 ;
        RECT 81.490 208.710 81.810 208.770 ;
        RECT 82.040 208.770 85.030 208.910 ;
        RECT 33.205 208.430 74.820 208.570 ;
        RECT 75.050 208.570 75.370 208.630 ;
        RECT 82.040 208.570 82.180 208.770 ;
        RECT 84.710 208.710 85.030 208.770 ;
        RECT 86.090 208.910 86.410 208.970 ;
        RECT 104.950 208.910 105.270 208.970 ;
        RECT 107.955 208.910 108.245 208.955 ;
        RECT 86.090 208.770 97.360 208.910 ;
        RECT 86.090 208.710 86.410 208.770 ;
        RECT 75.050 208.445 82.180 208.570 ;
        RECT 82.870 208.570 83.190 208.630 ;
        RECT 90.230 208.570 90.550 208.630 ;
        RECT 75.050 208.430 82.255 208.445 ;
        RECT 33.205 208.385 33.495 208.430 ;
        RECT 75.050 208.370 75.370 208.430 ;
        RECT 20.285 208.320 20.575 208.365 ;
        RECT 21.475 208.320 21.765 208.365 ;
        RECT 23.995 208.320 24.285 208.365 ;
        RECT 9.270 208.230 9.590 208.290 ;
        RECT 12.045 208.230 12.335 208.275 ;
        RECT 9.270 208.090 12.335 208.230 ;
        RECT 20.285 208.180 24.285 208.320 ;
        RECT 20.285 208.135 20.575 208.180 ;
        RECT 21.475 208.135 21.765 208.180 ;
        RECT 23.995 208.135 24.285 208.180 ;
        RECT 26.290 208.230 26.610 208.290 ;
        RECT 29.985 208.230 30.275 208.275 ;
        RECT 9.270 208.030 9.590 208.090 ;
        RECT 12.045 208.045 12.335 208.090 ;
        RECT 26.290 208.090 30.275 208.230 ;
        RECT 26.290 208.030 26.610 208.090 ;
        RECT 29.985 208.045 30.275 208.090 ;
        RECT 65.390 208.230 65.710 208.290 ;
        RECT 68.150 208.230 68.470 208.290 ;
        RECT 65.390 208.090 68.470 208.230 ;
        RECT 65.390 208.030 65.710 208.090 ;
        RECT 68.150 208.030 68.470 208.090 ;
        RECT 68.625 208.030 68.915 208.075 ;
        RECT 69.070 208.030 69.390 208.090 ;
        RECT 60.115 207.965 60.405 208.010 ;
        RECT 62.185 207.965 62.475 208.010 ;
        RECT 64.025 207.965 64.315 208.010 ;
        RECT 64.470 207.965 64.790 208.025 ;
        RECT 60.115 207.950 61.940 207.965 ;
        RECT 11.570 207.690 11.890 207.950 ;
        RECT 19.390 207.690 19.710 207.950 ;
        RECT 20.770 207.935 21.090 207.950 ;
        RECT 20.740 207.890 21.090 207.935 ;
        RECT 20.740 207.750 21.240 207.890 ;
        RECT 20.740 207.705 21.090 207.750 ;
        RECT 20.770 207.690 21.090 207.705 ;
        RECT 58.490 207.690 58.810 207.950 ;
        RECT 60.115 207.825 62.030 207.950 ;
        RECT 60.115 207.780 60.405 207.825 ;
        RECT 61.710 207.690 62.030 207.825 ;
        RECT 62.185 207.825 64.790 207.965 ;
        RECT 62.185 207.780 62.475 207.825 ;
        RECT 64.025 207.780 64.315 207.825 ;
        RECT 64.470 207.765 64.790 207.825 ;
        RECT 64.930 207.765 65.250 208.025 ;
        RECT 68.625 207.890 69.390 208.030 ;
        RECT 68.625 207.845 68.915 207.890 ;
        RECT 69.070 207.830 69.390 207.890 ;
        RECT 69.990 207.890 70.310 207.950 ;
        RECT 70.465 207.890 70.755 208.010 ;
        RECT 69.990 207.780 70.755 207.890 ;
        RECT 70.910 207.890 71.230 207.950 ;
        RECT 75.510 207.890 75.830 208.035 ;
        RECT 76.890 208.030 77.210 208.290 ;
        RECT 81.030 208.230 81.350 208.290 ;
        RECT 81.505 208.230 81.795 208.275 ;
        RECT 81.030 208.090 81.795 208.230 ;
        RECT 81.965 208.215 82.255 208.430 ;
        RECT 82.870 208.430 90.550 208.570 ;
        RECT 82.870 208.370 83.190 208.430 ;
        RECT 84.800 208.290 84.940 208.430 ;
        RECT 90.230 208.370 90.550 208.430 ;
        RECT 81.030 208.030 81.350 208.090 ;
        RECT 81.505 208.045 81.795 208.090 ;
        RECT 84.250 208.030 84.570 208.290 ;
        RECT 84.710 208.030 85.030 208.290 ;
        RECT 89.785 208.230 90.075 208.275 ;
        RECT 90.320 208.230 90.460 208.370 ;
        RECT 89.785 208.090 90.460 208.230 ;
        RECT 89.785 208.045 90.075 208.090 ;
        RECT 96.210 208.030 96.530 208.290 ;
        RECT 97.220 208.105 97.360 208.770 ;
        RECT 104.950 208.770 108.245 208.910 ;
        RECT 104.950 208.710 105.270 208.770 ;
        RECT 107.955 208.725 108.245 208.770 ;
        RECT 128.410 208.760 128.730 209.020 ;
        RECT 129.345 208.910 129.635 208.955 ;
        RECT 133.930 208.910 134.250 208.970 ;
        RECT 129.345 208.770 134.250 208.910 ;
        RECT 129.345 208.725 129.635 208.770 ;
        RECT 133.930 208.710 134.250 208.770 ;
        RECT 99.395 208.660 99.685 208.705 ;
        RECT 101.285 208.660 101.575 208.705 ;
        RECT 104.405 208.660 104.695 208.705 ;
        RECT 99.395 208.520 104.695 208.660 ;
        RECT 99.395 208.475 99.685 208.520 ;
        RECT 101.285 208.475 101.575 208.520 ;
        RECT 104.405 208.475 104.695 208.520 ;
        RECT 105.410 208.570 105.730 208.630 ;
        RECT 111.390 208.570 111.710 208.630 ;
        RECT 111.865 208.570 112.155 208.615 ;
        RECT 105.410 208.430 111.160 208.570 ;
        RECT 105.410 208.370 105.730 208.430 ;
        RECT 77.755 207.950 78.045 207.995 ;
        RECT 85.645 207.950 85.935 207.995 ;
        RECT 90.635 207.950 90.925 207.995 ;
        RECT 69.990 207.750 70.680 207.780 ;
        RECT 70.910 207.775 75.830 207.890 ;
        RECT 77.440 207.810 78.045 207.950 ;
        RECT 70.910 207.750 75.740 207.775 ;
        RECT 69.990 207.690 70.310 207.750 ;
        RECT 70.910 207.690 71.230 207.750 ;
        RECT 15.250 207.350 15.570 207.610 ;
        RECT 26.290 207.350 26.610 207.610 ;
        RECT 59.410 207.550 59.730 207.610 ;
        RECT 65.865 207.550 66.155 207.595 ;
        RECT 66.310 207.550 66.630 207.610 ;
        RECT 59.410 207.410 66.630 207.550 ;
        RECT 59.410 207.350 59.730 207.410 ;
        RECT 65.865 207.365 66.155 207.410 ;
        RECT 66.310 207.350 66.630 207.410 ;
        RECT 68.150 207.350 68.470 207.610 ;
        RECT 68.610 207.550 68.930 207.610 ;
        RECT 77.440 207.550 77.580 207.810 ;
        RECT 77.755 207.765 78.045 207.810 ;
        RECT 85.630 207.690 85.950 207.950 ;
        RECT 87.930 207.890 88.250 207.950 ;
        RECT 86.180 207.750 88.250 207.890 ;
        RECT 86.180 207.610 86.320 207.750 ;
        RECT 87.930 207.690 88.250 207.750 ;
        RECT 88.390 207.890 88.710 207.950 ;
        RECT 90.320 207.890 90.925 207.950 ;
        RECT 88.390 207.810 90.925 207.890 ;
        RECT 97.145 207.875 97.435 208.105 ;
        RECT 98.510 208.030 98.830 208.290 ;
        RECT 111.020 208.275 111.160 208.430 ;
        RECT 111.390 208.430 112.155 208.570 ;
        RECT 111.390 208.370 111.710 208.430 ;
        RECT 111.865 208.385 112.155 208.430 ;
        RECT 110.010 208.060 110.300 208.105 ;
        RECT 98.990 207.980 99.280 208.025 ;
        RECT 100.825 207.980 101.115 208.025 ;
        RECT 104.405 207.980 104.695 208.025 ;
        RECT 88.390 207.750 90.460 207.810 ;
        RECT 90.635 207.765 90.925 207.810 ;
        RECT 98.990 207.840 104.695 207.980 ;
        RECT 98.990 207.795 99.280 207.840 ;
        RECT 100.825 207.795 101.115 207.840 ;
        RECT 104.405 207.795 104.695 207.840 ;
        RECT 88.390 207.690 88.710 207.750 ;
        RECT 105.485 207.685 105.775 208.000 ;
        RECT 106.790 207.890 107.110 207.950 ;
        RECT 105.960 207.750 107.110 207.890 ;
        RECT 105.960 207.685 106.100 207.750 ;
        RECT 106.790 207.690 107.110 207.750 ;
        RECT 107.250 207.890 107.570 207.950 ;
        RECT 108.720 207.920 110.300 208.060 ;
        RECT 110.945 208.045 111.235 208.275 ;
        RECT 108.720 207.890 108.860 207.920 ;
        RECT 107.250 207.750 108.860 207.890 ;
        RECT 110.010 207.875 110.300 207.920 ;
        RECT 112.310 207.765 112.630 208.025 ;
        RECT 113.245 207.890 113.535 208.010 ;
        RECT 117.370 207.890 117.690 207.950 ;
        RECT 113.245 207.780 117.690 207.890 ;
        RECT 127.030 207.830 127.350 208.090 ;
        RECT 113.320 207.750 117.690 207.780 ;
        RECT 107.250 207.690 107.570 207.750 ;
        RECT 117.370 207.690 117.690 207.750 ;
        RECT 102.185 207.640 102.835 207.685 ;
        RECT 105.485 207.640 106.100 207.685 ;
        RECT 68.610 207.410 77.580 207.550 ;
        RECT 68.610 207.350 68.930 207.410 ;
        RECT 78.730 207.350 79.050 207.610 ;
        RECT 79.190 207.550 79.510 207.610 ;
        RECT 83.345 207.550 83.635 207.595 ;
        RECT 86.090 207.550 86.410 207.610 ;
        RECT 79.190 207.410 86.410 207.550 ;
        RECT 79.190 207.350 79.510 207.410 ;
        RECT 83.345 207.365 83.635 207.410 ;
        RECT 86.090 207.350 86.410 207.410 ;
        RECT 86.565 207.550 86.855 207.595 ;
        RECT 88.850 207.550 89.170 207.610 ;
        RECT 86.565 207.410 89.170 207.550 ;
        RECT 86.565 207.365 86.855 207.410 ;
        RECT 88.850 207.350 89.170 207.410 ;
        RECT 91.625 207.550 91.915 207.595 ;
        RECT 96.210 207.550 96.530 207.610 ;
        RECT 91.625 207.410 96.530 207.550 ;
        RECT 91.625 207.365 91.915 207.410 ;
        RECT 96.210 207.350 96.530 207.410 ;
        RECT 98.050 207.350 98.370 207.610 ;
        RECT 99.905 207.550 100.195 207.595 ;
        RECT 100.810 207.550 101.130 207.610 ;
        RECT 99.905 207.410 101.130 207.550 ;
        RECT 102.185 207.500 106.100 207.640 ;
        RECT 102.185 207.455 102.835 207.500 ;
        RECT 105.785 207.480 106.100 207.500 ;
        RECT 105.785 207.455 106.075 207.480 ;
        RECT 99.905 207.365 100.195 207.410 ;
        RECT 100.810 207.350 101.130 207.410 ;
        RECT 109.090 207.350 109.410 207.610 ;
        RECT 2.760 206.480 159.040 206.960 ;
        RECT 10.650 205.990 10.970 206.250 ;
        RECT 12.505 206.190 12.795 206.235 ;
        RECT 17.090 206.190 17.410 206.250 ;
        RECT 12.505 206.050 17.410 206.190 ;
        RECT 12.505 206.005 12.795 206.050 ;
        RECT 11.570 205.510 11.890 205.570 ;
        RECT 12.580 205.510 12.720 206.005 ;
        RECT 17.090 205.990 17.410 206.050 ;
        RECT 21.690 205.990 22.010 206.250 ;
        RECT 32.730 205.990 33.050 206.250 ;
        RECT 40.090 205.990 40.410 206.250 ;
        RECT 58.950 205.990 59.270 206.250 ;
        RECT 74.130 206.190 74.450 206.250 ;
        RECT 77.810 206.190 78.130 206.250 ;
        RECT 78.285 206.190 78.575 206.235 ;
        RECT 83.330 206.190 83.650 206.250 ;
        RECT 59.500 206.050 74.450 206.190 ;
        RECT 15.250 205.850 15.570 205.910 ;
        RECT 18.070 205.850 18.360 205.895 ;
        RECT 15.250 205.710 18.360 205.850 ;
        RECT 15.250 205.650 15.570 205.710 ;
        RECT 18.070 205.665 18.360 205.710 ;
        RECT 11.570 205.370 12.720 205.510 ;
        RECT 11.570 205.310 11.890 205.370 ;
        RECT 19.390 205.310 19.710 205.570 ;
        RECT 22.610 205.510 22.930 205.570 ;
        RECT 26.290 205.510 26.610 205.570 ;
        RECT 22.610 205.370 26.610 205.510 ;
        RECT 22.610 205.310 22.930 205.370 ;
        RECT 26.290 205.310 26.610 205.370 ;
        RECT 33.650 205.310 33.970 205.570 ;
        RECT 41.025 205.510 41.315 205.555 ;
        RECT 59.500 205.510 59.640 206.050 ;
        RECT 74.130 205.990 74.450 206.050 ;
        RECT 75.600 206.050 77.580 206.190 ;
        RECT 61.710 205.850 62.030 205.910 ;
        RECT 69.070 205.850 69.390 205.910 ;
        RECT 61.340 205.710 63.780 205.850 ;
        RECT 41.025 205.370 59.640 205.510 ;
        RECT 59.885 205.615 60.175 205.660 ;
        RECT 60.805 205.615 61.095 205.660 ;
        RECT 61.340 205.615 61.480 205.710 ;
        RECT 61.710 205.650 62.030 205.710 ;
        RECT 59.885 205.475 60.560 205.615 ;
        RECT 59.885 205.430 60.175 205.475 ;
        RECT 41.025 205.325 41.315 205.370 ;
        RECT 14.815 205.260 15.105 205.305 ;
        RECT 17.335 205.260 17.625 205.305 ;
        RECT 18.525 205.260 18.815 205.305 ;
        RECT 14.815 205.120 18.815 205.260 ;
        RECT 14.815 205.075 15.105 205.120 ;
        RECT 17.335 205.075 17.625 205.120 ;
        RECT 18.525 205.075 18.815 205.120 ;
        RECT 60.420 205.170 60.560 205.475 ;
        RECT 60.805 205.475 61.480 205.615 ;
        RECT 63.640 205.615 63.780 205.710 ;
        RECT 69.070 205.725 70.675 205.850 ;
        RECT 69.070 205.710 70.750 205.725 ;
        RECT 64.025 205.615 64.315 205.660 ;
        RECT 60.805 205.430 61.095 205.475 ;
        RECT 62.630 205.310 62.950 205.570 ;
        RECT 63.090 205.555 63.410 205.570 ;
        RECT 63.090 205.325 63.480 205.555 ;
        RECT 63.640 205.475 64.315 205.615 ;
        RECT 64.025 205.430 64.315 205.475 ;
        RECT 64.560 205.370 67.920 205.510 ;
        RECT 68.150 205.410 68.470 205.670 ;
        RECT 69.070 205.650 69.390 205.710 ;
        RECT 70.460 205.495 70.750 205.710 ;
        RECT 71.370 205.650 71.690 205.910 ;
        RECT 72.750 205.615 73.070 205.675 ;
        RECT 75.600 205.660 75.740 206.050 ;
        RECT 77.440 205.850 77.580 206.050 ;
        RECT 77.810 206.050 78.575 206.190 ;
        RECT 77.810 205.990 78.130 206.050 ;
        RECT 78.285 206.005 78.575 206.050 ;
        RECT 82.040 206.050 83.650 206.190 ;
        RECT 79.190 205.850 79.510 205.910 ;
        RECT 77.440 205.710 79.510 205.850 ;
        RECT 63.090 205.310 63.410 205.325 ;
        RECT 64.560 205.170 64.700 205.370 ;
        RECT 60.420 205.030 64.700 205.170 ;
        RECT 67.780 205.170 67.920 205.370 ;
        RECT 71.830 205.310 72.150 205.570 ;
        RECT 72.750 205.475 75.280 205.615 ;
        RECT 72.750 205.415 73.070 205.475 ;
        RECT 69.085 205.170 69.375 205.215 ;
        RECT 69.530 205.170 69.850 205.230 ;
        RECT 67.780 205.030 69.850 205.170 ;
        RECT 75.140 205.170 75.280 205.475 ;
        RECT 75.525 205.430 75.815 205.660 ;
        RECT 76.675 205.615 76.965 205.660 ;
        RECT 79.190 205.650 79.510 205.710 ;
        RECT 82.040 205.660 82.180 206.050 ;
        RECT 83.330 205.990 83.650 206.050 ;
        RECT 85.260 206.050 89.540 206.190 ;
        RECT 76.060 205.475 76.965 205.615 ;
        RECT 79.665 205.615 79.955 205.660 ;
        RECT 81.965 205.615 82.255 205.660 ;
        RECT 76.060 205.230 76.200 205.475 ;
        RECT 76.675 205.430 76.965 205.475 ;
        RECT 77.350 205.510 77.670 205.570 ;
        RECT 77.350 205.370 79.420 205.510 ;
        RECT 79.665 205.475 82.255 205.615 ;
        RECT 79.665 205.430 79.955 205.475 ;
        RECT 81.965 205.430 82.255 205.475 ;
        RECT 82.410 205.615 82.730 205.675 ;
        RECT 82.885 205.615 83.175 205.660 ;
        RECT 84.725 205.615 85.015 205.660 ;
        RECT 82.410 205.475 85.015 205.615 ;
        RECT 82.410 205.415 82.730 205.475 ;
        RECT 82.885 205.430 83.175 205.475 ;
        RECT 84.725 205.430 85.015 205.475 ;
        RECT 77.350 205.310 77.670 205.370 ;
        RECT 75.970 205.170 76.290 205.230 ;
        RECT 75.140 205.030 76.290 205.170 ;
        RECT 69.085 204.985 69.375 205.030 ;
        RECT 69.530 204.970 69.850 205.030 ;
        RECT 75.970 204.970 76.290 205.030 ;
        RECT 15.250 204.920 15.540 204.965 ;
        RECT 16.820 204.920 17.110 204.965 ;
        RECT 18.920 204.920 19.210 204.965 ;
        RECT 15.250 204.780 19.210 204.920 ;
        RECT 15.250 204.735 15.540 204.780 ;
        RECT 16.820 204.735 17.110 204.780 ;
        RECT 18.920 204.735 19.210 204.780 ;
        RECT 79.280 204.830 79.420 205.370 ;
        RECT 80.570 204.970 80.890 205.230 ;
        RECT 85.260 205.170 85.400 206.050 ;
        RECT 87.470 205.850 87.790 205.910 ;
        RECT 88.405 205.850 88.695 205.895 ;
        RECT 87.470 205.710 88.695 205.850 ;
        RECT 86.090 205.615 86.410 205.675 ;
        RECT 86.795 205.615 87.085 205.660 ;
        RECT 87.470 205.650 87.790 205.710 ;
        RECT 88.405 205.665 88.695 205.710 ;
        RECT 86.090 205.475 87.085 205.615 ;
        RECT 86.090 205.415 86.410 205.475 ;
        RECT 86.795 205.430 87.085 205.475 ;
        RECT 88.850 205.310 89.170 205.570 ;
        RECT 89.400 205.510 89.540 206.050 ;
        RECT 89.770 205.990 90.090 206.250 ;
        RECT 102.205 206.190 102.495 206.235 ;
        RECT 103.110 206.190 103.430 206.250 ;
        RECT 102.205 206.050 103.430 206.190 ;
        RECT 102.205 206.005 102.495 206.050 ;
        RECT 103.110 205.990 103.430 206.050 ;
        RECT 104.120 206.050 110.700 206.190 ;
        RECT 96.210 205.650 96.530 205.910 ;
        RECT 96.760 205.710 103.340 205.850 ;
        RECT 96.760 205.510 96.900 205.710 ;
        RECT 89.400 205.370 96.900 205.510 ;
        RECT 98.050 205.510 98.370 205.570 ;
        RECT 101.285 205.510 101.575 205.555 ;
        RECT 98.050 205.370 101.575 205.510 ;
        RECT 103.200 205.510 103.340 205.710 ;
        RECT 103.570 205.650 103.890 205.910 ;
        RECT 104.120 205.510 104.260 206.050 ;
        RECT 109.090 205.650 109.410 205.910 ;
        RECT 103.200 205.370 104.260 205.510 ;
        RECT 104.490 205.510 104.810 205.570 ;
        RECT 110.025 205.510 110.315 205.555 ;
        RECT 104.490 205.370 110.315 205.510 ;
        RECT 110.560 205.510 110.700 206.050 ;
        RECT 110.945 206.005 111.235 206.235 ;
        RECT 111.020 205.850 111.160 206.005 ;
        RECT 114.150 205.850 114.470 205.910 ;
        RECT 111.020 205.710 114.470 205.850 ;
        RECT 114.150 205.650 114.470 205.710 ;
        RECT 117.345 205.630 117.635 205.675 ;
        RECT 150.950 205.650 151.270 205.910 ;
        RECT 116.080 205.510 117.635 205.630 ;
        RECT 152.400 205.595 152.690 205.640 ;
        RECT 153.710 205.595 154.030 205.655 ;
        RECT 110.560 205.490 117.635 205.510 ;
        RECT 110.560 205.370 116.220 205.490 ;
        RECT 117.345 205.445 117.635 205.490 ;
        RECT 98.050 205.310 98.370 205.370 ;
        RECT 101.285 205.325 101.575 205.370 ;
        RECT 104.490 205.310 104.810 205.370 ;
        RECT 110.025 205.325 110.315 205.370 ;
        RECT 117.830 205.310 118.150 205.570 ;
        RECT 152.400 205.455 154.030 205.595 ;
        RECT 152.400 205.410 152.690 205.455 ;
        RECT 153.710 205.395 154.030 205.455 ;
        RECT 84.800 205.030 85.400 205.170 ;
        RECT 104.965 205.170 105.255 205.215 ;
        RECT 110.470 205.170 110.790 205.230 ;
        RECT 136.230 205.170 136.550 205.230 ;
        RECT 104.965 205.030 110.790 205.170 ;
        RECT 84.800 204.830 84.940 205.030 ;
        RECT 104.965 204.985 105.255 205.030 ;
        RECT 110.470 204.970 110.790 205.030 ;
        RECT 111.020 205.030 136.550 205.170 ;
        RECT 79.280 204.690 84.940 204.830 ;
        RECT 63.100 204.580 63.395 204.655 ;
        RECT 65.860 204.580 66.155 204.655 ;
        RECT 97.590 204.630 97.910 204.890 ;
        RECT 108.645 204.830 108.935 204.875 ;
        RECT 111.020 204.830 111.160 205.030 ;
        RECT 136.230 204.970 136.550 205.030 ;
        RECT 108.645 204.690 111.160 204.830 ;
        RECT 111.390 204.830 111.710 204.890 ;
        RECT 128.870 204.830 129.190 204.890 ;
        RECT 111.390 204.690 129.190 204.830 ;
        RECT 108.645 204.645 108.935 204.690 ;
        RECT 111.390 204.630 111.710 204.690 ;
        RECT 128.870 204.630 129.190 204.690 ;
        RECT 63.100 204.440 66.155 204.580 ;
        RECT 63.100 204.385 63.395 204.440 ;
        RECT 65.860 204.385 66.155 204.440 ;
        RECT 1.000 203.760 158.240 204.240 ;
        RECT 97.590 203.470 97.910 203.530 ;
        RECT 143.590 203.470 143.910 203.530 ;
        RECT 97.590 203.330 143.910 203.470 ;
        RECT 97.590 203.270 97.910 203.330 ;
        RECT 143.590 203.270 143.910 203.330 ;
        RECT 76.890 203.130 77.210 203.190 ;
        RECT 84.710 203.130 85.030 203.190 ;
        RECT 65.480 202.990 85.030 203.130 ;
        RECT 65.480 202.835 65.620 202.990 ;
        RECT 76.890 202.930 77.210 202.990 ;
        RECT 84.710 202.930 85.030 202.990 ;
        RECT 65.405 202.605 65.695 202.835 ;
        RECT 64.385 202.510 64.675 202.555 ;
        RECT 62.170 202.450 62.490 202.510 ;
        RECT 63.180 202.450 64.675 202.510 ;
        RECT 62.170 202.370 64.675 202.450 ;
        RECT 62.170 202.310 63.320 202.370 ;
        RECT 64.385 202.325 64.675 202.370 ;
        RECT 62.170 202.250 62.490 202.310 ;
        RECT 75.065 202.265 75.355 202.495 ;
        RECT 75.970 202.325 76.290 202.585 ;
        RECT 78.270 202.325 78.590 202.585 ;
        RECT 78.730 202.450 79.050 202.510 ;
        RECT 80.585 202.450 80.875 202.495 ;
        RECT 78.730 202.310 80.875 202.450 ;
        RECT 33.650 202.110 33.970 202.170 ;
        RECT 63.565 202.110 63.855 202.155 ;
        RECT 33.650 201.970 63.855 202.110 ;
        RECT 33.650 201.910 33.970 201.970 ;
        RECT 63.565 201.925 63.855 201.970 ;
        RECT 64.010 202.110 64.330 202.170 ;
        RECT 75.140 202.110 75.280 202.265 ;
        RECT 78.730 202.250 79.050 202.310 ;
        RECT 80.585 202.265 80.875 202.310 ;
        RECT 64.010 201.970 75.280 202.110 ;
        RECT 81.505 202.110 81.795 202.155 ;
        RECT 84.710 202.110 85.030 202.170 ;
        RECT 81.505 201.970 85.030 202.110 ;
        RECT 64.010 201.910 64.330 201.970 ;
        RECT 81.505 201.925 81.795 201.970 ;
        RECT 84.710 201.910 85.030 201.970 ;
        RECT 2.760 201.040 159.040 201.520 ;
        RECT 40.640 199.800 52.610 200.280 ;
        RECT 48.150 199.000 48.570 199.800 ;
        RECT 5.255 198.940 5.785 198.995 ;
        RECT 45.670 198.940 51.070 199.000 ;
        RECT 91.010 198.940 91.550 199.000 ;
        RECT 3.660 198.690 5.785 198.940 ;
        RECT 45.655 198.690 51.070 198.940 ;
        RECT 90.955 198.690 93.060 198.940 ;
        RECT 5.255 198.665 5.785 198.690 ;
        RECT 45.670 198.640 51.070 198.690 ;
        RECT 91.010 198.640 91.550 198.690 ;
        RECT 48.150 197.800 48.570 198.640 ;
        RECT 157.490 197.800 158.960 198.820 ;
        RECT 1.100 197.410 158.960 197.800 ;
        RECT 10.250 158.495 10.600 166.485 ;
        RECT 11.600 165.585 19.700 165.885 ;
        RECT 11.320 163.160 11.550 165.405 ;
        RECT 11.275 161.760 11.735 163.160 ;
        RECT 11.320 159.405 11.550 161.760 ;
        RECT 11.960 160.960 12.190 165.405 ;
        RECT 12.600 163.160 12.830 165.405 ;
        RECT 12.550 161.760 13.010 163.160 ;
        RECT 11.925 159.560 12.385 160.960 ;
        RECT 11.960 159.405 12.190 159.560 ;
        RECT 12.600 159.405 12.830 161.760 ;
        RECT 13.240 160.960 13.470 165.405 ;
        RECT 13.880 163.160 14.110 165.405 ;
        RECT 13.825 161.760 14.285 163.160 ;
        RECT 13.215 159.560 13.675 160.960 ;
        RECT 13.240 159.405 13.470 159.560 ;
        RECT 13.880 159.405 14.110 161.760 ;
        RECT 14.520 160.960 14.750 165.405 ;
        RECT 15.160 163.160 15.390 165.405 ;
        RECT 15.100 161.760 15.560 163.160 ;
        RECT 14.490 159.560 14.950 160.960 ;
        RECT 14.520 159.405 14.750 159.560 ;
        RECT 15.160 159.405 15.390 161.760 ;
        RECT 15.800 160.960 16.030 165.405 ;
        RECT 16.440 163.160 16.670 165.405 ;
        RECT 16.375 161.760 16.835 163.160 ;
        RECT 15.765 159.560 16.225 160.960 ;
        RECT 15.800 159.405 16.030 159.560 ;
        RECT 16.440 159.405 16.670 161.760 ;
        RECT 17.080 160.960 17.310 165.405 ;
        RECT 17.720 163.160 17.950 165.405 ;
        RECT 17.650 161.760 18.110 163.160 ;
        RECT 17.040 159.560 17.500 160.960 ;
        RECT 17.080 159.405 17.310 159.560 ;
        RECT 17.720 159.405 17.950 161.760 ;
        RECT 18.360 160.960 18.590 165.405 ;
        RECT 19.300 164.410 19.700 165.585 ;
        RECT 25.350 164.410 25.700 164.460 ;
        RECT 19.300 164.110 25.700 164.410 ;
        RECT 18.315 159.560 18.775 160.960 ;
        RECT 18.360 159.405 18.590 159.560 ;
        RECT 19.300 159.210 19.700 164.110 ;
        RECT 25.350 164.060 25.700 164.110 ;
        RECT 21.550 163.510 25.700 163.810 ;
        RECT 21.280 163.160 21.510 163.360 ;
        RECT 21.225 161.760 21.685 163.160 ;
        RECT 21.280 159.360 21.510 161.760 ;
        RECT 21.920 160.960 22.150 163.360 ;
        RECT 22.560 163.160 22.790 163.360 ;
        RECT 22.500 161.760 22.960 163.160 ;
        RECT 21.890 159.560 22.350 160.960 ;
        RECT 21.920 159.360 22.150 159.560 ;
        RECT 22.560 159.360 22.790 161.760 ;
        RECT 23.200 160.960 23.430 163.360 ;
        RECT 23.840 163.160 24.070 163.360 ;
        RECT 23.775 161.760 24.235 163.160 ;
        RECT 23.165 159.560 23.625 160.960 ;
        RECT 23.200 159.360 23.430 159.560 ;
        RECT 23.840 159.360 24.070 161.760 ;
        RECT 24.480 160.960 24.710 163.360 ;
        RECT 25.430 162.760 25.700 163.510 ;
        RECT 25.350 162.360 25.700 162.760 ;
        RECT 24.450 159.560 24.810 160.960 ;
        RECT 24.480 159.360 24.710 159.560 ;
        RECT 25.430 159.210 25.700 162.360 ;
        RECT 11.600 158.910 19.700 159.210 ;
        RECT 8.050 157.430 17.300 158.495 ;
        RECT 17.920 158.010 18.150 158.100 ;
        RECT 18.360 158.010 18.590 158.100 ;
        RECT 19.300 158.010 19.700 158.910 ;
        RECT 20.160 158.910 25.700 159.210 ;
        RECT 17.815 157.660 18.175 158.010 ;
        RECT 18.340 157.660 18.700 158.010 ;
        RECT 19.250 157.660 19.750 158.010 ;
        RECT 17.920 157.100 18.150 157.660 ;
        RECT 18.360 157.100 18.590 157.660 ;
        RECT 19.300 157.610 19.700 157.660 ;
        RECT 16.600 156.910 17.050 156.960 ;
        RECT 20.160 156.910 20.560 158.910 ;
        RECT 25.850 158.760 26.200 166.480 ;
        RECT 22.670 158.560 26.200 158.760 ;
        RECT 21.280 158.010 21.510 158.070 ;
        RECT 21.720 158.010 21.950 158.070 ;
        RECT 21.165 157.660 21.525 158.010 ;
        RECT 21.690 157.660 22.050 158.010 ;
        RECT 22.670 157.660 23.200 158.560 ;
        RECT 25.100 158.495 26.200 158.560 ;
        RECT 23.920 158.010 24.150 158.060 ;
        RECT 23.775 157.660 24.150 158.010 ;
        RECT 21.280 157.070 21.510 157.660 ;
        RECT 21.720 157.070 21.950 157.660 ;
        RECT 23.920 157.060 24.150 157.660 ;
        RECT 24.360 158.010 24.590 158.060 ;
        RECT 24.360 157.660 24.740 158.010 ;
        RECT 24.360 157.060 24.590 157.660 ;
        RECT 25.100 157.430 26.335 158.495 ;
        RECT 133.790 158.485 134.140 166.475 ;
        RECT 134.290 165.875 134.640 165.925 ;
        RECT 134.290 165.575 143.240 165.875 ;
        RECT 134.860 163.150 135.090 165.395 ;
        RECT 134.815 161.750 135.275 163.150 ;
        RECT 134.860 159.395 135.090 161.750 ;
        RECT 135.500 160.950 135.730 165.395 ;
        RECT 136.140 163.150 136.370 165.395 ;
        RECT 136.090 161.750 136.550 163.150 ;
        RECT 135.465 159.550 135.925 160.950 ;
        RECT 135.500 159.395 135.730 159.550 ;
        RECT 136.140 159.395 136.370 161.750 ;
        RECT 136.780 160.950 137.010 165.395 ;
        RECT 137.420 163.150 137.650 165.395 ;
        RECT 137.365 161.750 137.825 163.150 ;
        RECT 136.755 159.550 137.215 160.950 ;
        RECT 136.780 159.395 137.010 159.550 ;
        RECT 137.420 159.395 137.650 161.750 ;
        RECT 138.060 160.950 138.290 165.395 ;
        RECT 138.700 163.150 138.930 165.395 ;
        RECT 138.640 161.750 139.100 163.150 ;
        RECT 138.030 159.550 138.490 160.950 ;
        RECT 138.060 159.395 138.290 159.550 ;
        RECT 138.700 159.395 138.930 161.750 ;
        RECT 139.340 160.950 139.570 165.395 ;
        RECT 139.980 163.150 140.210 165.395 ;
        RECT 139.915 161.750 140.375 163.150 ;
        RECT 139.305 159.550 139.765 160.950 ;
        RECT 139.340 159.395 139.570 159.550 ;
        RECT 139.980 159.395 140.210 161.750 ;
        RECT 140.620 160.950 140.850 165.395 ;
        RECT 141.260 163.150 141.490 165.395 ;
        RECT 141.190 161.750 141.650 163.150 ;
        RECT 140.580 159.550 141.040 160.950 ;
        RECT 140.620 159.395 140.850 159.550 ;
        RECT 141.260 159.395 141.490 161.750 ;
        RECT 141.900 160.950 142.130 165.395 ;
        RECT 141.855 159.550 142.315 160.950 ;
        RECT 141.900 159.395 142.130 159.550 ;
        RECT 142.840 159.200 143.240 165.575 ;
        RECT 145.090 163.500 149.240 163.800 ;
        RECT 144.820 163.150 145.050 163.350 ;
        RECT 144.765 161.750 145.225 163.150 ;
        RECT 144.820 159.350 145.050 161.750 ;
        RECT 145.460 160.950 145.690 163.350 ;
        RECT 146.100 163.150 146.330 163.350 ;
        RECT 146.040 161.750 146.500 163.150 ;
        RECT 145.430 159.550 145.890 160.950 ;
        RECT 145.460 159.350 145.690 159.550 ;
        RECT 146.100 159.350 146.330 161.750 ;
        RECT 146.740 160.950 146.970 163.350 ;
        RECT 147.380 163.150 147.610 163.350 ;
        RECT 147.315 161.750 147.775 163.150 ;
        RECT 146.705 159.550 147.165 160.950 ;
        RECT 146.740 159.350 146.970 159.550 ;
        RECT 147.380 159.350 147.610 161.750 ;
        RECT 148.020 160.950 148.250 163.350 ;
        RECT 147.990 159.550 148.350 160.950 ;
        RECT 148.020 159.350 148.250 159.550 ;
        RECT 148.970 159.200 149.240 163.500 ;
        RECT 135.140 158.900 143.240 159.200 ;
        RECT 145.090 158.900 149.240 159.200 ;
        RECT 16.600 156.680 21.760 156.910 ;
        RECT 16.600 156.660 21.735 156.680 ;
        RECT 16.600 156.610 17.050 156.660 ;
        RECT 24.025 156.595 24.475 156.915 ;
        RECT 10.250 148.495 10.600 156.485 ;
        RECT 11.600 155.585 19.700 155.885 ;
        RECT 11.320 153.160 11.550 155.405 ;
        RECT 11.275 151.760 11.735 153.160 ;
        RECT 11.320 149.405 11.550 151.760 ;
        RECT 11.960 150.960 12.190 155.405 ;
        RECT 12.600 153.160 12.830 155.405 ;
        RECT 12.550 151.760 13.010 153.160 ;
        RECT 11.925 149.560 12.385 150.960 ;
        RECT 11.960 149.405 12.190 149.560 ;
        RECT 12.600 149.405 12.830 151.760 ;
        RECT 13.240 150.960 13.470 155.405 ;
        RECT 13.880 153.160 14.110 155.405 ;
        RECT 13.825 151.760 14.285 153.160 ;
        RECT 13.215 149.560 13.675 150.960 ;
        RECT 13.240 149.405 13.470 149.560 ;
        RECT 13.880 149.405 14.110 151.760 ;
        RECT 14.520 150.960 14.750 155.405 ;
        RECT 15.160 153.160 15.390 155.405 ;
        RECT 15.100 151.760 15.560 153.160 ;
        RECT 14.490 149.560 14.950 150.960 ;
        RECT 14.520 149.405 14.750 149.560 ;
        RECT 15.160 149.405 15.390 151.760 ;
        RECT 15.800 150.960 16.030 155.405 ;
        RECT 16.440 153.160 16.670 155.405 ;
        RECT 16.375 151.760 16.835 153.160 ;
        RECT 15.765 149.560 16.225 150.960 ;
        RECT 15.800 149.405 16.030 149.560 ;
        RECT 16.440 149.405 16.670 151.760 ;
        RECT 17.080 150.960 17.310 155.405 ;
        RECT 17.720 153.160 17.950 155.405 ;
        RECT 17.650 151.760 18.110 153.160 ;
        RECT 17.040 149.560 17.500 150.960 ;
        RECT 17.080 149.405 17.310 149.560 ;
        RECT 17.720 149.405 17.950 151.760 ;
        RECT 18.360 150.960 18.590 155.405 ;
        RECT 19.300 154.410 19.700 155.585 ;
        RECT 25.350 154.410 25.700 154.460 ;
        RECT 19.300 154.110 25.700 154.410 ;
        RECT 18.315 149.560 18.775 150.960 ;
        RECT 18.360 149.405 18.590 149.560 ;
        RECT 19.300 149.210 19.700 154.110 ;
        RECT 25.350 154.060 25.700 154.110 ;
        RECT 21.550 153.510 25.700 153.810 ;
        RECT 21.280 153.160 21.510 153.360 ;
        RECT 21.225 151.760 21.685 153.160 ;
        RECT 21.280 149.360 21.510 151.760 ;
        RECT 21.920 150.960 22.150 153.360 ;
        RECT 22.560 153.160 22.790 153.360 ;
        RECT 22.500 151.760 22.960 153.160 ;
        RECT 21.890 149.560 22.350 150.960 ;
        RECT 21.920 149.360 22.150 149.560 ;
        RECT 22.560 149.360 22.790 151.760 ;
        RECT 23.200 150.960 23.430 153.360 ;
        RECT 23.840 153.160 24.070 153.360 ;
        RECT 23.775 151.760 24.235 153.160 ;
        RECT 23.165 149.560 23.625 150.960 ;
        RECT 23.200 149.360 23.430 149.560 ;
        RECT 23.840 149.360 24.070 151.760 ;
        RECT 24.480 150.960 24.710 153.360 ;
        RECT 25.430 152.760 25.700 153.510 ;
        RECT 25.350 152.360 25.700 152.760 ;
        RECT 24.450 149.560 24.810 150.960 ;
        RECT 24.480 149.360 24.710 149.560 ;
        RECT 25.430 149.210 25.700 152.360 ;
        RECT 11.600 148.910 19.700 149.210 ;
        RECT 8.050 147.430 17.300 148.495 ;
        RECT 17.920 148.010 18.150 148.100 ;
        RECT 18.360 148.010 18.590 148.100 ;
        RECT 19.300 148.010 19.700 148.910 ;
        RECT 20.160 148.910 25.700 149.210 ;
        RECT 17.815 147.660 18.175 148.010 ;
        RECT 18.340 147.660 18.700 148.010 ;
        RECT 19.250 147.660 19.750 148.010 ;
        RECT 17.920 147.100 18.150 147.660 ;
        RECT 18.360 147.100 18.590 147.660 ;
        RECT 19.300 147.610 19.700 147.660 ;
        RECT 16.600 146.910 17.050 146.960 ;
        RECT 20.160 146.910 20.560 148.910 ;
        RECT 25.850 148.760 26.200 157.430 ;
        RECT 133.655 157.420 140.840 158.485 ;
        RECT 141.460 158.000 141.690 158.090 ;
        RECT 141.900 158.000 142.130 158.090 ;
        RECT 142.840 158.000 143.240 158.900 ;
        RECT 144.820 158.000 145.050 158.060 ;
        RECT 145.260 158.000 145.490 158.060 ;
        RECT 141.355 157.650 141.715 158.000 ;
        RECT 141.880 157.650 142.240 158.000 ;
        RECT 142.790 157.650 143.290 158.000 ;
        RECT 144.705 157.650 145.065 158.000 ;
        RECT 145.230 157.650 145.590 158.000 ;
        RECT 141.460 157.090 141.690 157.650 ;
        RECT 141.900 157.090 142.130 157.650 ;
        RECT 142.840 157.600 143.240 157.650 ;
        RECT 144.820 157.060 145.050 157.650 ;
        RECT 145.260 157.060 145.490 157.650 ;
        RECT 146.390 156.955 146.690 158.900 ;
        RECT 149.390 158.485 149.740 166.475 ;
        RECT 146.840 157.420 151.990 158.485 ;
        RECT 139.690 156.900 140.090 156.950 ;
        RECT 146.335 156.900 146.745 156.955 ;
        RECT 139.690 156.650 146.745 156.900 ;
        RECT 139.690 156.600 140.090 156.650 ;
        RECT 146.335 156.595 146.745 156.650 ;
        RECT 22.670 148.560 26.200 148.760 ;
        RECT 21.280 148.010 21.510 148.070 ;
        RECT 21.720 148.010 21.950 148.070 ;
        RECT 21.165 147.660 21.525 148.010 ;
        RECT 21.690 147.660 22.050 148.010 ;
        RECT 22.670 147.660 23.200 148.560 ;
        RECT 25.100 148.495 26.200 148.560 ;
        RECT 23.920 148.010 24.150 148.060 ;
        RECT 23.775 147.660 24.150 148.010 ;
        RECT 21.280 147.070 21.510 147.660 ;
        RECT 21.720 147.070 21.950 147.660 ;
        RECT 23.920 147.060 24.150 147.660 ;
        RECT 24.360 148.010 24.590 148.060 ;
        RECT 24.360 147.660 24.740 148.010 ;
        RECT 24.360 147.060 24.590 147.660 ;
        RECT 25.100 147.430 26.335 148.495 ;
        RECT 133.790 148.485 134.140 156.475 ;
        RECT 134.290 155.875 134.640 155.925 ;
        RECT 134.290 155.575 143.240 155.875 ;
        RECT 134.860 153.150 135.090 155.395 ;
        RECT 134.815 151.750 135.275 153.150 ;
        RECT 134.860 149.395 135.090 151.750 ;
        RECT 135.500 150.950 135.730 155.395 ;
        RECT 136.140 153.150 136.370 155.395 ;
        RECT 136.090 151.750 136.550 153.150 ;
        RECT 135.465 149.550 135.925 150.950 ;
        RECT 135.500 149.395 135.730 149.550 ;
        RECT 136.140 149.395 136.370 151.750 ;
        RECT 136.780 150.950 137.010 155.395 ;
        RECT 137.420 153.150 137.650 155.395 ;
        RECT 137.365 151.750 137.825 153.150 ;
        RECT 136.755 149.550 137.215 150.950 ;
        RECT 136.780 149.395 137.010 149.550 ;
        RECT 137.420 149.395 137.650 151.750 ;
        RECT 138.060 150.950 138.290 155.395 ;
        RECT 138.700 153.150 138.930 155.395 ;
        RECT 138.640 151.750 139.100 153.150 ;
        RECT 138.030 149.550 138.490 150.950 ;
        RECT 138.060 149.395 138.290 149.550 ;
        RECT 138.700 149.395 138.930 151.750 ;
        RECT 139.340 150.950 139.570 155.395 ;
        RECT 139.980 153.150 140.210 155.395 ;
        RECT 139.915 151.750 140.375 153.150 ;
        RECT 139.305 149.550 139.765 150.950 ;
        RECT 139.340 149.395 139.570 149.550 ;
        RECT 139.980 149.395 140.210 151.750 ;
        RECT 140.620 150.950 140.850 155.395 ;
        RECT 141.260 153.150 141.490 155.395 ;
        RECT 141.190 151.750 141.650 153.150 ;
        RECT 140.580 149.550 141.040 150.950 ;
        RECT 140.620 149.395 140.850 149.550 ;
        RECT 141.260 149.395 141.490 151.750 ;
        RECT 141.900 150.950 142.130 155.395 ;
        RECT 141.855 149.550 142.315 150.950 ;
        RECT 141.900 149.395 142.130 149.550 ;
        RECT 142.840 149.200 143.240 155.575 ;
        RECT 145.090 153.500 149.240 153.800 ;
        RECT 144.820 153.150 145.050 153.350 ;
        RECT 144.765 151.750 145.225 153.150 ;
        RECT 144.820 149.350 145.050 151.750 ;
        RECT 145.460 150.950 145.690 153.350 ;
        RECT 146.100 153.150 146.330 153.350 ;
        RECT 146.040 151.750 146.500 153.150 ;
        RECT 145.430 149.550 145.890 150.950 ;
        RECT 145.460 149.350 145.690 149.550 ;
        RECT 146.100 149.350 146.330 151.750 ;
        RECT 146.740 150.950 146.970 153.350 ;
        RECT 147.380 153.150 147.610 153.350 ;
        RECT 147.315 151.750 147.775 153.150 ;
        RECT 146.705 149.550 147.165 150.950 ;
        RECT 146.740 149.350 146.970 149.550 ;
        RECT 147.380 149.350 147.610 151.750 ;
        RECT 148.020 150.950 148.250 153.350 ;
        RECT 147.990 149.550 148.350 150.950 ;
        RECT 148.020 149.350 148.250 149.550 ;
        RECT 148.970 149.200 149.240 153.500 ;
        RECT 135.140 148.900 143.240 149.200 ;
        RECT 145.090 148.900 149.240 149.200 ;
        RECT 16.600 146.680 21.760 146.910 ;
        RECT 16.600 146.660 21.735 146.680 ;
        RECT 16.600 146.610 17.050 146.660 ;
        RECT 24.025 146.595 24.475 146.915 ;
        RECT 10.250 138.495 10.600 146.485 ;
        RECT 11.600 145.585 19.700 145.885 ;
        RECT 11.320 143.160 11.550 145.405 ;
        RECT 11.275 141.760 11.735 143.160 ;
        RECT 11.320 139.405 11.550 141.760 ;
        RECT 11.960 140.960 12.190 145.405 ;
        RECT 12.600 143.160 12.830 145.405 ;
        RECT 12.550 141.760 13.010 143.160 ;
        RECT 11.925 139.560 12.385 140.960 ;
        RECT 11.960 139.405 12.190 139.560 ;
        RECT 12.600 139.405 12.830 141.760 ;
        RECT 13.240 140.960 13.470 145.405 ;
        RECT 13.880 143.160 14.110 145.405 ;
        RECT 13.825 141.760 14.285 143.160 ;
        RECT 13.215 139.560 13.675 140.960 ;
        RECT 13.240 139.405 13.470 139.560 ;
        RECT 13.880 139.405 14.110 141.760 ;
        RECT 14.520 140.960 14.750 145.405 ;
        RECT 15.160 143.160 15.390 145.405 ;
        RECT 15.100 141.760 15.560 143.160 ;
        RECT 14.490 139.560 14.950 140.960 ;
        RECT 14.520 139.405 14.750 139.560 ;
        RECT 15.160 139.405 15.390 141.760 ;
        RECT 15.800 140.960 16.030 145.405 ;
        RECT 16.440 143.160 16.670 145.405 ;
        RECT 16.375 141.760 16.835 143.160 ;
        RECT 15.765 139.560 16.225 140.960 ;
        RECT 15.800 139.405 16.030 139.560 ;
        RECT 16.440 139.405 16.670 141.760 ;
        RECT 17.080 140.960 17.310 145.405 ;
        RECT 17.720 143.160 17.950 145.405 ;
        RECT 17.650 141.760 18.110 143.160 ;
        RECT 17.040 139.560 17.500 140.960 ;
        RECT 17.080 139.405 17.310 139.560 ;
        RECT 17.720 139.405 17.950 141.760 ;
        RECT 18.360 140.960 18.590 145.405 ;
        RECT 19.300 144.410 19.700 145.585 ;
        RECT 25.350 144.410 25.700 144.460 ;
        RECT 19.300 144.110 25.700 144.410 ;
        RECT 18.315 139.560 18.775 140.960 ;
        RECT 18.360 139.405 18.590 139.560 ;
        RECT 19.300 139.210 19.700 144.110 ;
        RECT 25.350 144.060 25.700 144.110 ;
        RECT 21.550 143.510 25.700 143.810 ;
        RECT 21.280 143.160 21.510 143.360 ;
        RECT 21.225 141.760 21.685 143.160 ;
        RECT 21.280 139.360 21.510 141.760 ;
        RECT 21.920 140.960 22.150 143.360 ;
        RECT 22.560 143.160 22.790 143.360 ;
        RECT 22.500 141.760 22.960 143.160 ;
        RECT 21.890 139.560 22.350 140.960 ;
        RECT 21.920 139.360 22.150 139.560 ;
        RECT 22.560 139.360 22.790 141.760 ;
        RECT 23.200 140.960 23.430 143.360 ;
        RECT 23.840 143.160 24.070 143.360 ;
        RECT 23.775 141.760 24.235 143.160 ;
        RECT 23.165 139.560 23.625 140.960 ;
        RECT 23.200 139.360 23.430 139.560 ;
        RECT 23.840 139.360 24.070 141.760 ;
        RECT 24.480 140.960 24.710 143.360 ;
        RECT 25.430 142.760 25.700 143.510 ;
        RECT 25.350 142.360 25.700 142.760 ;
        RECT 24.450 139.560 24.810 140.960 ;
        RECT 24.480 139.360 24.710 139.560 ;
        RECT 25.430 139.210 25.700 142.360 ;
        RECT 11.600 138.910 19.700 139.210 ;
        RECT 8.050 137.430 17.300 138.495 ;
        RECT 17.920 138.010 18.150 138.100 ;
        RECT 18.360 138.010 18.590 138.100 ;
        RECT 19.300 138.010 19.700 138.910 ;
        RECT 20.160 138.910 25.700 139.210 ;
        RECT 17.815 137.660 18.175 138.010 ;
        RECT 18.340 137.660 18.700 138.010 ;
        RECT 19.250 137.660 19.750 138.010 ;
        RECT 17.920 137.100 18.150 137.660 ;
        RECT 18.360 137.100 18.590 137.660 ;
        RECT 19.300 137.610 19.700 137.660 ;
        RECT 16.600 136.910 17.050 136.960 ;
        RECT 20.160 136.910 20.560 138.910 ;
        RECT 25.850 138.760 26.200 147.430 ;
        RECT 133.655 147.420 140.840 148.485 ;
        RECT 141.460 148.000 141.690 148.090 ;
        RECT 141.900 148.000 142.130 148.090 ;
        RECT 142.840 148.000 143.240 148.900 ;
        RECT 144.820 148.000 145.050 148.060 ;
        RECT 145.260 148.000 145.490 148.060 ;
        RECT 141.355 147.650 141.715 148.000 ;
        RECT 141.880 147.650 142.240 148.000 ;
        RECT 142.790 147.650 143.290 148.000 ;
        RECT 144.705 147.650 145.065 148.000 ;
        RECT 145.230 147.650 145.590 148.000 ;
        RECT 141.460 147.090 141.690 147.650 ;
        RECT 141.900 147.090 142.130 147.650 ;
        RECT 142.840 147.600 143.240 147.650 ;
        RECT 144.820 147.060 145.050 147.650 ;
        RECT 145.260 147.060 145.490 147.650 ;
        RECT 146.390 146.955 146.690 148.900 ;
        RECT 149.390 148.485 149.740 156.475 ;
        RECT 146.840 147.420 151.990 148.485 ;
        RECT 139.690 146.900 140.090 146.950 ;
        RECT 146.335 146.900 146.745 146.955 ;
        RECT 139.690 146.650 146.745 146.900 ;
        RECT 139.690 146.600 140.090 146.650 ;
        RECT 146.335 146.595 146.745 146.650 ;
        RECT 22.670 138.560 26.200 138.760 ;
        RECT 21.280 138.010 21.510 138.070 ;
        RECT 21.720 138.010 21.950 138.070 ;
        RECT 21.165 137.660 21.525 138.010 ;
        RECT 21.690 137.660 22.050 138.010 ;
        RECT 22.670 137.660 23.200 138.560 ;
        RECT 25.100 138.495 26.200 138.560 ;
        RECT 23.920 138.010 24.150 138.060 ;
        RECT 23.775 137.660 24.150 138.010 ;
        RECT 21.280 137.070 21.510 137.660 ;
        RECT 21.720 137.070 21.950 137.660 ;
        RECT 23.920 137.060 24.150 137.660 ;
        RECT 24.360 138.010 24.590 138.060 ;
        RECT 24.360 137.660 24.740 138.010 ;
        RECT 24.360 137.060 24.590 137.660 ;
        RECT 25.100 137.430 26.335 138.495 ;
        RECT 133.790 138.485 134.140 146.475 ;
        RECT 134.290 145.875 134.640 145.925 ;
        RECT 134.290 145.575 143.240 145.875 ;
        RECT 134.860 143.150 135.090 145.395 ;
        RECT 134.815 141.750 135.275 143.150 ;
        RECT 134.860 139.395 135.090 141.750 ;
        RECT 135.500 140.950 135.730 145.395 ;
        RECT 136.140 143.150 136.370 145.395 ;
        RECT 136.090 141.750 136.550 143.150 ;
        RECT 135.465 139.550 135.925 140.950 ;
        RECT 135.500 139.395 135.730 139.550 ;
        RECT 136.140 139.395 136.370 141.750 ;
        RECT 136.780 140.950 137.010 145.395 ;
        RECT 137.420 143.150 137.650 145.395 ;
        RECT 137.365 141.750 137.825 143.150 ;
        RECT 136.755 139.550 137.215 140.950 ;
        RECT 136.780 139.395 137.010 139.550 ;
        RECT 137.420 139.395 137.650 141.750 ;
        RECT 138.060 140.950 138.290 145.395 ;
        RECT 138.700 143.150 138.930 145.395 ;
        RECT 138.640 141.750 139.100 143.150 ;
        RECT 138.030 139.550 138.490 140.950 ;
        RECT 138.060 139.395 138.290 139.550 ;
        RECT 138.700 139.395 138.930 141.750 ;
        RECT 139.340 140.950 139.570 145.395 ;
        RECT 139.980 143.150 140.210 145.395 ;
        RECT 139.915 141.750 140.375 143.150 ;
        RECT 139.305 139.550 139.765 140.950 ;
        RECT 139.340 139.395 139.570 139.550 ;
        RECT 139.980 139.395 140.210 141.750 ;
        RECT 140.620 140.950 140.850 145.395 ;
        RECT 141.260 143.150 141.490 145.395 ;
        RECT 141.190 141.750 141.650 143.150 ;
        RECT 140.580 139.550 141.040 140.950 ;
        RECT 140.620 139.395 140.850 139.550 ;
        RECT 141.260 139.395 141.490 141.750 ;
        RECT 141.900 140.950 142.130 145.395 ;
        RECT 141.855 139.550 142.315 140.950 ;
        RECT 141.900 139.395 142.130 139.550 ;
        RECT 142.840 139.200 143.240 145.575 ;
        RECT 145.090 143.500 149.240 143.800 ;
        RECT 144.820 143.150 145.050 143.350 ;
        RECT 144.765 141.750 145.225 143.150 ;
        RECT 144.820 139.350 145.050 141.750 ;
        RECT 145.460 140.950 145.690 143.350 ;
        RECT 146.100 143.150 146.330 143.350 ;
        RECT 146.040 141.750 146.500 143.150 ;
        RECT 145.430 139.550 145.890 140.950 ;
        RECT 145.460 139.350 145.690 139.550 ;
        RECT 146.100 139.350 146.330 141.750 ;
        RECT 146.740 140.950 146.970 143.350 ;
        RECT 147.380 143.150 147.610 143.350 ;
        RECT 147.315 141.750 147.775 143.150 ;
        RECT 146.705 139.550 147.165 140.950 ;
        RECT 146.740 139.350 146.970 139.550 ;
        RECT 147.380 139.350 147.610 141.750 ;
        RECT 148.020 140.950 148.250 143.350 ;
        RECT 147.990 139.550 148.350 140.950 ;
        RECT 148.020 139.350 148.250 139.550 ;
        RECT 148.970 139.200 149.240 143.500 ;
        RECT 135.140 138.900 143.240 139.200 ;
        RECT 145.090 138.900 149.240 139.200 ;
        RECT 16.600 136.680 21.760 136.910 ;
        RECT 16.600 136.660 21.735 136.680 ;
        RECT 16.600 136.610 17.050 136.660 ;
        RECT 24.025 136.595 24.475 136.915 ;
        RECT 10.250 128.495 10.600 136.485 ;
        RECT 11.600 135.585 19.700 135.885 ;
        RECT 11.320 133.160 11.550 135.405 ;
        RECT 11.275 131.760 11.735 133.160 ;
        RECT 11.320 129.405 11.550 131.760 ;
        RECT 11.960 130.960 12.190 135.405 ;
        RECT 12.600 133.160 12.830 135.405 ;
        RECT 12.550 131.760 13.010 133.160 ;
        RECT 11.925 129.560 12.385 130.960 ;
        RECT 11.960 129.405 12.190 129.560 ;
        RECT 12.600 129.405 12.830 131.760 ;
        RECT 13.240 130.960 13.470 135.405 ;
        RECT 13.880 133.160 14.110 135.405 ;
        RECT 13.825 131.760 14.285 133.160 ;
        RECT 13.215 129.560 13.675 130.960 ;
        RECT 13.240 129.405 13.470 129.560 ;
        RECT 13.880 129.405 14.110 131.760 ;
        RECT 14.520 130.960 14.750 135.405 ;
        RECT 15.160 133.160 15.390 135.405 ;
        RECT 15.100 131.760 15.560 133.160 ;
        RECT 14.490 129.560 14.950 130.960 ;
        RECT 14.520 129.405 14.750 129.560 ;
        RECT 15.160 129.405 15.390 131.760 ;
        RECT 15.800 130.960 16.030 135.405 ;
        RECT 16.440 133.160 16.670 135.405 ;
        RECT 16.375 131.760 16.835 133.160 ;
        RECT 15.765 129.560 16.225 130.960 ;
        RECT 15.800 129.405 16.030 129.560 ;
        RECT 16.440 129.405 16.670 131.760 ;
        RECT 17.080 130.960 17.310 135.405 ;
        RECT 17.720 133.160 17.950 135.405 ;
        RECT 17.650 131.760 18.110 133.160 ;
        RECT 17.040 129.560 17.500 130.960 ;
        RECT 17.080 129.405 17.310 129.560 ;
        RECT 17.720 129.405 17.950 131.760 ;
        RECT 18.360 130.960 18.590 135.405 ;
        RECT 19.300 134.410 19.700 135.585 ;
        RECT 25.350 134.410 25.700 134.460 ;
        RECT 19.300 134.110 25.700 134.410 ;
        RECT 18.315 129.560 18.775 130.960 ;
        RECT 18.360 129.405 18.590 129.560 ;
        RECT 19.300 129.210 19.700 134.110 ;
        RECT 25.350 134.060 25.700 134.110 ;
        RECT 21.550 133.510 25.700 133.810 ;
        RECT 21.280 133.160 21.510 133.360 ;
        RECT 21.225 131.760 21.685 133.160 ;
        RECT 21.280 129.360 21.510 131.760 ;
        RECT 21.920 130.960 22.150 133.360 ;
        RECT 22.560 133.160 22.790 133.360 ;
        RECT 22.500 131.760 22.960 133.160 ;
        RECT 21.890 129.560 22.350 130.960 ;
        RECT 21.920 129.360 22.150 129.560 ;
        RECT 22.560 129.360 22.790 131.760 ;
        RECT 23.200 130.960 23.430 133.360 ;
        RECT 23.840 133.160 24.070 133.360 ;
        RECT 23.775 131.760 24.235 133.160 ;
        RECT 23.165 129.560 23.625 130.960 ;
        RECT 23.200 129.360 23.430 129.560 ;
        RECT 23.840 129.360 24.070 131.760 ;
        RECT 24.480 130.960 24.710 133.360 ;
        RECT 25.430 132.760 25.700 133.510 ;
        RECT 25.350 132.360 25.700 132.760 ;
        RECT 24.450 129.560 24.810 130.960 ;
        RECT 24.480 129.360 24.710 129.560 ;
        RECT 25.430 129.210 25.700 132.360 ;
        RECT 11.600 128.910 19.700 129.210 ;
        RECT 8.050 127.430 17.300 128.495 ;
        RECT 17.920 128.010 18.150 128.100 ;
        RECT 18.360 128.010 18.590 128.100 ;
        RECT 19.300 128.010 19.700 128.910 ;
        RECT 20.160 128.910 25.700 129.210 ;
        RECT 17.815 127.660 18.175 128.010 ;
        RECT 18.340 127.660 18.700 128.010 ;
        RECT 19.250 127.660 19.750 128.010 ;
        RECT 17.920 127.100 18.150 127.660 ;
        RECT 18.360 127.100 18.590 127.660 ;
        RECT 19.300 127.610 19.700 127.660 ;
        RECT 16.600 126.910 17.050 126.960 ;
        RECT 20.160 126.910 20.560 128.910 ;
        RECT 25.850 128.760 26.200 137.430 ;
        RECT 133.655 137.420 140.840 138.485 ;
        RECT 141.460 138.000 141.690 138.090 ;
        RECT 141.900 138.000 142.130 138.090 ;
        RECT 142.840 138.000 143.240 138.900 ;
        RECT 144.820 138.000 145.050 138.060 ;
        RECT 145.260 138.000 145.490 138.060 ;
        RECT 141.355 137.650 141.715 138.000 ;
        RECT 141.880 137.650 142.240 138.000 ;
        RECT 142.790 137.650 143.290 138.000 ;
        RECT 144.705 137.650 145.065 138.000 ;
        RECT 145.230 137.650 145.590 138.000 ;
        RECT 141.460 137.090 141.690 137.650 ;
        RECT 141.900 137.090 142.130 137.650 ;
        RECT 142.840 137.600 143.240 137.650 ;
        RECT 144.820 137.060 145.050 137.650 ;
        RECT 145.260 137.060 145.490 137.650 ;
        RECT 146.390 136.955 146.690 138.900 ;
        RECT 149.390 138.485 149.740 146.475 ;
        RECT 146.840 137.420 151.990 138.485 ;
        RECT 139.690 136.900 140.090 136.950 ;
        RECT 146.335 136.900 146.745 136.955 ;
        RECT 139.690 136.650 146.745 136.900 ;
        RECT 139.690 136.600 140.090 136.650 ;
        RECT 146.335 136.595 146.745 136.650 ;
        RECT 22.670 128.560 26.200 128.760 ;
        RECT 21.280 128.010 21.510 128.070 ;
        RECT 21.720 128.010 21.950 128.070 ;
        RECT 21.165 127.660 21.525 128.010 ;
        RECT 21.690 127.660 22.050 128.010 ;
        RECT 22.670 127.660 23.200 128.560 ;
        RECT 25.100 128.495 26.200 128.560 ;
        RECT 23.920 128.010 24.150 128.060 ;
        RECT 23.775 127.660 24.150 128.010 ;
        RECT 21.280 127.070 21.510 127.660 ;
        RECT 21.720 127.070 21.950 127.660 ;
        RECT 23.920 127.060 24.150 127.660 ;
        RECT 24.360 128.010 24.590 128.060 ;
        RECT 24.360 127.660 24.740 128.010 ;
        RECT 24.360 127.060 24.590 127.660 ;
        RECT 25.100 127.430 26.335 128.495 ;
        RECT 133.790 128.485 134.140 136.475 ;
        RECT 134.290 135.875 134.640 135.925 ;
        RECT 134.290 135.575 143.240 135.875 ;
        RECT 134.860 133.150 135.090 135.395 ;
        RECT 134.815 131.750 135.275 133.150 ;
        RECT 134.860 129.395 135.090 131.750 ;
        RECT 135.500 130.950 135.730 135.395 ;
        RECT 136.140 133.150 136.370 135.395 ;
        RECT 136.090 131.750 136.550 133.150 ;
        RECT 135.465 129.550 135.925 130.950 ;
        RECT 135.500 129.395 135.730 129.550 ;
        RECT 136.140 129.395 136.370 131.750 ;
        RECT 136.780 130.950 137.010 135.395 ;
        RECT 137.420 133.150 137.650 135.395 ;
        RECT 137.365 131.750 137.825 133.150 ;
        RECT 136.755 129.550 137.215 130.950 ;
        RECT 136.780 129.395 137.010 129.550 ;
        RECT 137.420 129.395 137.650 131.750 ;
        RECT 138.060 130.950 138.290 135.395 ;
        RECT 138.700 133.150 138.930 135.395 ;
        RECT 138.640 131.750 139.100 133.150 ;
        RECT 138.030 129.550 138.490 130.950 ;
        RECT 138.060 129.395 138.290 129.550 ;
        RECT 138.700 129.395 138.930 131.750 ;
        RECT 139.340 130.950 139.570 135.395 ;
        RECT 139.980 133.150 140.210 135.395 ;
        RECT 139.915 131.750 140.375 133.150 ;
        RECT 139.305 129.550 139.765 130.950 ;
        RECT 139.340 129.395 139.570 129.550 ;
        RECT 139.980 129.395 140.210 131.750 ;
        RECT 140.620 130.950 140.850 135.395 ;
        RECT 141.260 133.150 141.490 135.395 ;
        RECT 141.190 131.750 141.650 133.150 ;
        RECT 140.580 129.550 141.040 130.950 ;
        RECT 140.620 129.395 140.850 129.550 ;
        RECT 141.260 129.395 141.490 131.750 ;
        RECT 141.900 130.950 142.130 135.395 ;
        RECT 141.855 129.550 142.315 130.950 ;
        RECT 141.900 129.395 142.130 129.550 ;
        RECT 142.840 129.200 143.240 135.575 ;
        RECT 145.090 133.500 149.240 133.800 ;
        RECT 144.820 133.150 145.050 133.350 ;
        RECT 144.765 131.750 145.225 133.150 ;
        RECT 144.820 129.350 145.050 131.750 ;
        RECT 145.460 130.950 145.690 133.350 ;
        RECT 146.100 133.150 146.330 133.350 ;
        RECT 146.040 131.750 146.500 133.150 ;
        RECT 145.430 129.550 145.890 130.950 ;
        RECT 145.460 129.350 145.690 129.550 ;
        RECT 146.100 129.350 146.330 131.750 ;
        RECT 146.740 130.950 146.970 133.350 ;
        RECT 147.380 133.150 147.610 133.350 ;
        RECT 147.315 131.750 147.775 133.150 ;
        RECT 146.705 129.550 147.165 130.950 ;
        RECT 146.740 129.350 146.970 129.550 ;
        RECT 147.380 129.350 147.610 131.750 ;
        RECT 148.020 130.950 148.250 133.350 ;
        RECT 147.990 129.550 148.350 130.950 ;
        RECT 148.020 129.350 148.250 129.550 ;
        RECT 148.970 129.200 149.240 133.500 ;
        RECT 135.140 128.900 143.240 129.200 ;
        RECT 145.090 128.900 149.240 129.200 ;
        RECT 16.600 126.680 21.760 126.910 ;
        RECT 16.600 126.660 21.735 126.680 ;
        RECT 16.600 126.610 17.050 126.660 ;
        RECT 24.025 126.595 24.475 126.915 ;
        RECT 10.250 118.495 10.600 126.485 ;
        RECT 11.600 125.585 19.700 125.885 ;
        RECT 11.320 123.160 11.550 125.405 ;
        RECT 11.275 121.760 11.735 123.160 ;
        RECT 11.320 119.405 11.550 121.760 ;
        RECT 11.960 120.960 12.190 125.405 ;
        RECT 12.600 123.160 12.830 125.405 ;
        RECT 12.550 121.760 13.010 123.160 ;
        RECT 11.925 119.560 12.385 120.960 ;
        RECT 11.960 119.405 12.190 119.560 ;
        RECT 12.600 119.405 12.830 121.760 ;
        RECT 13.240 120.960 13.470 125.405 ;
        RECT 13.880 123.160 14.110 125.405 ;
        RECT 13.825 121.760 14.285 123.160 ;
        RECT 13.215 119.560 13.675 120.960 ;
        RECT 13.240 119.405 13.470 119.560 ;
        RECT 13.880 119.405 14.110 121.760 ;
        RECT 14.520 120.960 14.750 125.405 ;
        RECT 15.160 123.160 15.390 125.405 ;
        RECT 15.100 121.760 15.560 123.160 ;
        RECT 14.490 119.560 14.950 120.960 ;
        RECT 14.520 119.405 14.750 119.560 ;
        RECT 15.160 119.405 15.390 121.760 ;
        RECT 15.800 120.960 16.030 125.405 ;
        RECT 16.440 123.160 16.670 125.405 ;
        RECT 16.375 121.760 16.835 123.160 ;
        RECT 15.765 119.560 16.225 120.960 ;
        RECT 15.800 119.405 16.030 119.560 ;
        RECT 16.440 119.405 16.670 121.760 ;
        RECT 17.080 120.960 17.310 125.405 ;
        RECT 17.720 123.160 17.950 125.405 ;
        RECT 17.650 121.760 18.110 123.160 ;
        RECT 17.040 119.560 17.500 120.960 ;
        RECT 17.080 119.405 17.310 119.560 ;
        RECT 17.720 119.405 17.950 121.760 ;
        RECT 18.360 120.960 18.590 125.405 ;
        RECT 19.300 124.410 19.700 125.585 ;
        RECT 25.350 124.410 25.700 124.460 ;
        RECT 19.300 124.110 25.700 124.410 ;
        RECT 18.315 119.560 18.775 120.960 ;
        RECT 18.360 119.405 18.590 119.560 ;
        RECT 19.300 119.210 19.700 124.110 ;
        RECT 25.350 124.060 25.700 124.110 ;
        RECT 21.550 123.510 25.700 123.810 ;
        RECT 21.280 123.160 21.510 123.360 ;
        RECT 21.225 121.760 21.685 123.160 ;
        RECT 21.280 119.360 21.510 121.760 ;
        RECT 21.920 120.960 22.150 123.360 ;
        RECT 22.560 123.160 22.790 123.360 ;
        RECT 22.500 121.760 22.960 123.160 ;
        RECT 21.890 119.560 22.350 120.960 ;
        RECT 21.920 119.360 22.150 119.560 ;
        RECT 22.560 119.360 22.790 121.760 ;
        RECT 23.200 120.960 23.430 123.360 ;
        RECT 23.840 123.160 24.070 123.360 ;
        RECT 23.775 121.760 24.235 123.160 ;
        RECT 23.165 119.560 23.625 120.960 ;
        RECT 23.200 119.360 23.430 119.560 ;
        RECT 23.840 119.360 24.070 121.760 ;
        RECT 24.480 120.960 24.710 123.360 ;
        RECT 25.430 122.760 25.700 123.510 ;
        RECT 25.350 122.360 25.700 122.760 ;
        RECT 24.450 119.560 24.810 120.960 ;
        RECT 24.480 119.360 24.710 119.560 ;
        RECT 25.430 119.210 25.700 122.360 ;
        RECT 11.600 118.910 19.700 119.210 ;
        RECT 8.050 117.430 17.300 118.495 ;
        RECT 17.920 118.010 18.150 118.100 ;
        RECT 18.360 118.010 18.590 118.100 ;
        RECT 19.300 118.010 19.700 118.910 ;
        RECT 20.160 118.910 25.700 119.210 ;
        RECT 17.815 117.660 18.175 118.010 ;
        RECT 18.340 117.660 18.700 118.010 ;
        RECT 19.250 117.660 19.750 118.010 ;
        RECT 17.920 117.100 18.150 117.660 ;
        RECT 18.360 117.100 18.590 117.660 ;
        RECT 19.300 117.610 19.700 117.660 ;
        RECT 16.600 116.910 17.050 116.960 ;
        RECT 20.160 116.910 20.560 118.910 ;
        RECT 25.850 118.760 26.200 127.430 ;
        RECT 133.655 127.420 140.840 128.485 ;
        RECT 141.460 128.000 141.690 128.090 ;
        RECT 141.900 128.000 142.130 128.090 ;
        RECT 142.840 128.000 143.240 128.900 ;
        RECT 144.820 128.000 145.050 128.060 ;
        RECT 145.260 128.000 145.490 128.060 ;
        RECT 141.355 127.650 141.715 128.000 ;
        RECT 141.880 127.650 142.240 128.000 ;
        RECT 142.790 127.650 143.290 128.000 ;
        RECT 144.705 127.650 145.065 128.000 ;
        RECT 145.230 127.650 145.590 128.000 ;
        RECT 141.460 127.090 141.690 127.650 ;
        RECT 141.900 127.090 142.130 127.650 ;
        RECT 142.840 127.600 143.240 127.650 ;
        RECT 144.820 127.060 145.050 127.650 ;
        RECT 145.260 127.060 145.490 127.650 ;
        RECT 146.390 126.955 146.690 128.900 ;
        RECT 149.390 128.485 149.740 136.475 ;
        RECT 146.840 127.420 151.990 128.485 ;
        RECT 139.690 126.900 140.090 126.950 ;
        RECT 146.335 126.900 146.745 126.955 ;
        RECT 139.690 126.650 146.745 126.900 ;
        RECT 139.690 126.600 140.090 126.650 ;
        RECT 146.335 126.595 146.745 126.650 ;
        RECT 22.670 118.560 26.200 118.760 ;
        RECT 21.280 118.010 21.510 118.070 ;
        RECT 21.720 118.010 21.950 118.070 ;
        RECT 21.165 117.660 21.525 118.010 ;
        RECT 21.690 117.660 22.050 118.010 ;
        RECT 22.670 117.660 23.200 118.560 ;
        RECT 25.100 118.495 26.200 118.560 ;
        RECT 23.920 118.010 24.150 118.060 ;
        RECT 23.775 117.660 24.150 118.010 ;
        RECT 21.280 117.070 21.510 117.660 ;
        RECT 21.720 117.070 21.950 117.660 ;
        RECT 23.920 117.060 24.150 117.660 ;
        RECT 24.360 118.010 24.590 118.060 ;
        RECT 24.360 117.660 24.740 118.010 ;
        RECT 24.360 117.060 24.590 117.660 ;
        RECT 25.100 117.430 26.335 118.495 ;
        RECT 133.790 118.485 134.140 126.475 ;
        RECT 134.290 125.875 134.640 125.925 ;
        RECT 134.290 125.575 143.240 125.875 ;
        RECT 134.860 123.150 135.090 125.395 ;
        RECT 134.815 121.750 135.275 123.150 ;
        RECT 134.860 119.395 135.090 121.750 ;
        RECT 135.500 120.950 135.730 125.395 ;
        RECT 136.140 123.150 136.370 125.395 ;
        RECT 136.090 121.750 136.550 123.150 ;
        RECT 135.465 119.550 135.925 120.950 ;
        RECT 135.500 119.395 135.730 119.550 ;
        RECT 136.140 119.395 136.370 121.750 ;
        RECT 136.780 120.950 137.010 125.395 ;
        RECT 137.420 123.150 137.650 125.395 ;
        RECT 137.365 121.750 137.825 123.150 ;
        RECT 136.755 119.550 137.215 120.950 ;
        RECT 136.780 119.395 137.010 119.550 ;
        RECT 137.420 119.395 137.650 121.750 ;
        RECT 138.060 120.950 138.290 125.395 ;
        RECT 138.700 123.150 138.930 125.395 ;
        RECT 138.640 121.750 139.100 123.150 ;
        RECT 138.030 119.550 138.490 120.950 ;
        RECT 138.060 119.395 138.290 119.550 ;
        RECT 138.700 119.395 138.930 121.750 ;
        RECT 139.340 120.950 139.570 125.395 ;
        RECT 139.980 123.150 140.210 125.395 ;
        RECT 139.915 121.750 140.375 123.150 ;
        RECT 139.305 119.550 139.765 120.950 ;
        RECT 139.340 119.395 139.570 119.550 ;
        RECT 139.980 119.395 140.210 121.750 ;
        RECT 140.620 120.950 140.850 125.395 ;
        RECT 141.260 123.150 141.490 125.395 ;
        RECT 141.190 121.750 141.650 123.150 ;
        RECT 140.580 119.550 141.040 120.950 ;
        RECT 140.620 119.395 140.850 119.550 ;
        RECT 141.260 119.395 141.490 121.750 ;
        RECT 141.900 120.950 142.130 125.395 ;
        RECT 141.855 119.550 142.315 120.950 ;
        RECT 141.900 119.395 142.130 119.550 ;
        RECT 142.840 119.200 143.240 125.575 ;
        RECT 145.090 123.500 149.240 123.800 ;
        RECT 144.820 123.150 145.050 123.350 ;
        RECT 144.765 121.750 145.225 123.150 ;
        RECT 144.820 119.350 145.050 121.750 ;
        RECT 145.460 120.950 145.690 123.350 ;
        RECT 146.100 123.150 146.330 123.350 ;
        RECT 146.040 121.750 146.500 123.150 ;
        RECT 145.430 119.550 145.890 120.950 ;
        RECT 145.460 119.350 145.690 119.550 ;
        RECT 146.100 119.350 146.330 121.750 ;
        RECT 146.740 120.950 146.970 123.350 ;
        RECT 147.380 123.150 147.610 123.350 ;
        RECT 147.315 121.750 147.775 123.150 ;
        RECT 146.705 119.550 147.165 120.950 ;
        RECT 146.740 119.350 146.970 119.550 ;
        RECT 147.380 119.350 147.610 121.750 ;
        RECT 148.020 120.950 148.250 123.350 ;
        RECT 147.990 119.550 148.350 120.950 ;
        RECT 148.020 119.350 148.250 119.550 ;
        RECT 148.970 119.200 149.240 123.500 ;
        RECT 135.140 118.900 143.240 119.200 ;
        RECT 145.090 118.900 149.240 119.200 ;
        RECT 16.600 116.680 21.760 116.910 ;
        RECT 16.600 116.660 21.735 116.680 ;
        RECT 16.600 116.610 17.050 116.660 ;
        RECT 24.025 116.595 24.475 116.915 ;
        RECT 10.250 108.495 10.600 116.485 ;
        RECT 11.600 115.585 19.700 115.885 ;
        RECT 11.320 113.160 11.550 115.405 ;
        RECT 11.275 111.760 11.735 113.160 ;
        RECT 11.320 109.405 11.550 111.760 ;
        RECT 11.960 110.960 12.190 115.405 ;
        RECT 12.600 113.160 12.830 115.405 ;
        RECT 12.550 111.760 13.010 113.160 ;
        RECT 11.925 109.560 12.385 110.960 ;
        RECT 11.960 109.405 12.190 109.560 ;
        RECT 12.600 109.405 12.830 111.760 ;
        RECT 13.240 110.960 13.470 115.405 ;
        RECT 13.880 113.160 14.110 115.405 ;
        RECT 13.825 111.760 14.285 113.160 ;
        RECT 13.215 109.560 13.675 110.960 ;
        RECT 13.240 109.405 13.470 109.560 ;
        RECT 13.880 109.405 14.110 111.760 ;
        RECT 14.520 110.960 14.750 115.405 ;
        RECT 15.160 113.160 15.390 115.405 ;
        RECT 15.100 111.760 15.560 113.160 ;
        RECT 14.490 109.560 14.950 110.960 ;
        RECT 14.520 109.405 14.750 109.560 ;
        RECT 15.160 109.405 15.390 111.760 ;
        RECT 15.800 110.960 16.030 115.405 ;
        RECT 16.440 113.160 16.670 115.405 ;
        RECT 16.375 111.760 16.835 113.160 ;
        RECT 15.765 109.560 16.225 110.960 ;
        RECT 15.800 109.405 16.030 109.560 ;
        RECT 16.440 109.405 16.670 111.760 ;
        RECT 17.080 110.960 17.310 115.405 ;
        RECT 17.720 113.160 17.950 115.405 ;
        RECT 17.650 111.760 18.110 113.160 ;
        RECT 17.040 109.560 17.500 110.960 ;
        RECT 17.080 109.405 17.310 109.560 ;
        RECT 17.720 109.405 17.950 111.760 ;
        RECT 18.360 110.960 18.590 115.405 ;
        RECT 19.300 114.410 19.700 115.585 ;
        RECT 25.350 114.410 25.700 114.460 ;
        RECT 19.300 114.110 25.700 114.410 ;
        RECT 18.315 109.560 18.775 110.960 ;
        RECT 18.360 109.405 18.590 109.560 ;
        RECT 19.300 109.210 19.700 114.110 ;
        RECT 25.350 114.060 25.700 114.110 ;
        RECT 21.550 113.510 25.700 113.810 ;
        RECT 21.280 113.160 21.510 113.360 ;
        RECT 21.225 111.760 21.685 113.160 ;
        RECT 21.280 109.360 21.510 111.760 ;
        RECT 21.920 110.960 22.150 113.360 ;
        RECT 22.560 113.160 22.790 113.360 ;
        RECT 22.500 111.760 22.960 113.160 ;
        RECT 21.890 109.560 22.350 110.960 ;
        RECT 21.920 109.360 22.150 109.560 ;
        RECT 22.560 109.360 22.790 111.760 ;
        RECT 23.200 110.960 23.430 113.360 ;
        RECT 23.840 113.160 24.070 113.360 ;
        RECT 23.775 111.760 24.235 113.160 ;
        RECT 23.165 109.560 23.625 110.960 ;
        RECT 23.200 109.360 23.430 109.560 ;
        RECT 23.840 109.360 24.070 111.760 ;
        RECT 24.480 110.960 24.710 113.360 ;
        RECT 25.430 112.760 25.700 113.510 ;
        RECT 25.350 112.360 25.700 112.760 ;
        RECT 24.450 109.560 24.810 110.960 ;
        RECT 24.480 109.360 24.710 109.560 ;
        RECT 25.430 109.210 25.700 112.360 ;
        RECT 11.600 108.910 19.700 109.210 ;
        RECT 8.050 107.430 17.300 108.495 ;
        RECT 17.920 108.010 18.150 108.100 ;
        RECT 18.360 108.010 18.590 108.100 ;
        RECT 19.300 108.010 19.700 108.910 ;
        RECT 20.160 108.910 25.700 109.210 ;
        RECT 17.815 107.660 18.175 108.010 ;
        RECT 18.340 107.660 18.700 108.010 ;
        RECT 19.250 107.660 19.750 108.010 ;
        RECT 17.920 107.100 18.150 107.660 ;
        RECT 18.360 107.100 18.590 107.660 ;
        RECT 19.300 107.610 19.700 107.660 ;
        RECT 16.600 106.910 17.050 106.960 ;
        RECT 20.160 106.910 20.560 108.910 ;
        RECT 25.850 108.760 26.200 117.430 ;
        RECT 133.655 117.420 140.840 118.485 ;
        RECT 141.460 118.000 141.690 118.090 ;
        RECT 141.900 118.000 142.130 118.090 ;
        RECT 142.840 118.000 143.240 118.900 ;
        RECT 144.820 118.000 145.050 118.060 ;
        RECT 145.260 118.000 145.490 118.060 ;
        RECT 141.355 117.650 141.715 118.000 ;
        RECT 141.880 117.650 142.240 118.000 ;
        RECT 142.790 117.650 143.290 118.000 ;
        RECT 144.705 117.650 145.065 118.000 ;
        RECT 145.230 117.650 145.590 118.000 ;
        RECT 141.460 117.090 141.690 117.650 ;
        RECT 141.900 117.090 142.130 117.650 ;
        RECT 142.840 117.600 143.240 117.650 ;
        RECT 144.820 117.060 145.050 117.650 ;
        RECT 145.260 117.060 145.490 117.650 ;
        RECT 146.390 116.955 146.690 118.900 ;
        RECT 149.390 118.485 149.740 126.475 ;
        RECT 146.840 117.420 151.990 118.485 ;
        RECT 139.690 116.900 140.090 116.950 ;
        RECT 146.335 116.900 146.745 116.955 ;
        RECT 139.690 116.650 146.745 116.900 ;
        RECT 139.690 116.600 140.090 116.650 ;
        RECT 146.335 116.595 146.745 116.650 ;
        RECT 22.670 108.560 26.200 108.760 ;
        RECT 21.280 108.010 21.510 108.070 ;
        RECT 21.720 108.010 21.950 108.070 ;
        RECT 21.165 107.660 21.525 108.010 ;
        RECT 21.690 107.660 22.050 108.010 ;
        RECT 22.670 107.660 23.200 108.560 ;
        RECT 25.100 108.495 26.200 108.560 ;
        RECT 23.920 108.010 24.150 108.060 ;
        RECT 23.775 107.660 24.150 108.010 ;
        RECT 21.280 107.070 21.510 107.660 ;
        RECT 21.720 107.070 21.950 107.660 ;
        RECT 23.920 107.060 24.150 107.660 ;
        RECT 24.360 108.010 24.590 108.060 ;
        RECT 24.360 107.660 24.740 108.010 ;
        RECT 24.360 107.060 24.590 107.660 ;
        RECT 25.100 107.430 26.335 108.495 ;
        RECT 133.790 108.485 134.140 116.475 ;
        RECT 134.290 115.875 134.640 115.925 ;
        RECT 134.290 115.575 143.240 115.875 ;
        RECT 134.860 113.150 135.090 115.395 ;
        RECT 134.815 111.750 135.275 113.150 ;
        RECT 134.860 109.395 135.090 111.750 ;
        RECT 135.500 110.950 135.730 115.395 ;
        RECT 136.140 113.150 136.370 115.395 ;
        RECT 136.090 111.750 136.550 113.150 ;
        RECT 135.465 109.550 135.925 110.950 ;
        RECT 135.500 109.395 135.730 109.550 ;
        RECT 136.140 109.395 136.370 111.750 ;
        RECT 136.780 110.950 137.010 115.395 ;
        RECT 137.420 113.150 137.650 115.395 ;
        RECT 137.365 111.750 137.825 113.150 ;
        RECT 136.755 109.550 137.215 110.950 ;
        RECT 136.780 109.395 137.010 109.550 ;
        RECT 137.420 109.395 137.650 111.750 ;
        RECT 138.060 110.950 138.290 115.395 ;
        RECT 138.700 113.150 138.930 115.395 ;
        RECT 138.640 111.750 139.100 113.150 ;
        RECT 138.030 109.550 138.490 110.950 ;
        RECT 138.060 109.395 138.290 109.550 ;
        RECT 138.700 109.395 138.930 111.750 ;
        RECT 139.340 110.950 139.570 115.395 ;
        RECT 139.980 113.150 140.210 115.395 ;
        RECT 139.915 111.750 140.375 113.150 ;
        RECT 139.305 109.550 139.765 110.950 ;
        RECT 139.340 109.395 139.570 109.550 ;
        RECT 139.980 109.395 140.210 111.750 ;
        RECT 140.620 110.950 140.850 115.395 ;
        RECT 141.260 113.150 141.490 115.395 ;
        RECT 141.190 111.750 141.650 113.150 ;
        RECT 140.580 109.550 141.040 110.950 ;
        RECT 140.620 109.395 140.850 109.550 ;
        RECT 141.260 109.395 141.490 111.750 ;
        RECT 141.900 110.950 142.130 115.395 ;
        RECT 141.855 109.550 142.315 110.950 ;
        RECT 141.900 109.395 142.130 109.550 ;
        RECT 142.840 109.200 143.240 115.575 ;
        RECT 145.090 113.500 149.240 113.800 ;
        RECT 144.820 113.150 145.050 113.350 ;
        RECT 144.765 111.750 145.225 113.150 ;
        RECT 144.820 109.350 145.050 111.750 ;
        RECT 145.460 110.950 145.690 113.350 ;
        RECT 146.100 113.150 146.330 113.350 ;
        RECT 146.040 111.750 146.500 113.150 ;
        RECT 145.430 109.550 145.890 110.950 ;
        RECT 145.460 109.350 145.690 109.550 ;
        RECT 146.100 109.350 146.330 111.750 ;
        RECT 146.740 110.950 146.970 113.350 ;
        RECT 147.380 113.150 147.610 113.350 ;
        RECT 147.315 111.750 147.775 113.150 ;
        RECT 146.705 109.550 147.165 110.950 ;
        RECT 146.740 109.350 146.970 109.550 ;
        RECT 147.380 109.350 147.610 111.750 ;
        RECT 148.020 110.950 148.250 113.350 ;
        RECT 147.990 109.550 148.350 110.950 ;
        RECT 148.020 109.350 148.250 109.550 ;
        RECT 148.970 109.200 149.240 113.500 ;
        RECT 135.140 108.900 143.240 109.200 ;
        RECT 145.090 108.900 149.240 109.200 ;
        RECT 16.600 106.680 21.760 106.910 ;
        RECT 16.600 106.660 21.735 106.680 ;
        RECT 16.600 106.610 17.050 106.660 ;
        RECT 24.025 106.595 24.475 106.915 ;
        RECT 10.250 98.495 10.600 106.485 ;
        RECT 11.600 105.585 19.700 105.885 ;
        RECT 11.320 103.160 11.550 105.405 ;
        RECT 11.275 101.760 11.735 103.160 ;
        RECT 11.320 99.405 11.550 101.760 ;
        RECT 11.960 100.960 12.190 105.405 ;
        RECT 12.600 103.160 12.830 105.405 ;
        RECT 12.550 101.760 13.010 103.160 ;
        RECT 11.925 99.560 12.385 100.960 ;
        RECT 11.960 99.405 12.190 99.560 ;
        RECT 12.600 99.405 12.830 101.760 ;
        RECT 13.240 100.960 13.470 105.405 ;
        RECT 13.880 103.160 14.110 105.405 ;
        RECT 13.825 101.760 14.285 103.160 ;
        RECT 13.215 99.560 13.675 100.960 ;
        RECT 13.240 99.405 13.470 99.560 ;
        RECT 13.880 99.405 14.110 101.760 ;
        RECT 14.520 100.960 14.750 105.405 ;
        RECT 15.160 103.160 15.390 105.405 ;
        RECT 15.100 101.760 15.560 103.160 ;
        RECT 14.490 99.560 14.950 100.960 ;
        RECT 14.520 99.405 14.750 99.560 ;
        RECT 15.160 99.405 15.390 101.760 ;
        RECT 15.800 100.960 16.030 105.405 ;
        RECT 16.440 103.160 16.670 105.405 ;
        RECT 16.375 101.760 16.835 103.160 ;
        RECT 15.765 99.560 16.225 100.960 ;
        RECT 15.800 99.405 16.030 99.560 ;
        RECT 16.440 99.405 16.670 101.760 ;
        RECT 17.080 100.960 17.310 105.405 ;
        RECT 17.720 103.160 17.950 105.405 ;
        RECT 17.650 101.760 18.110 103.160 ;
        RECT 17.040 99.560 17.500 100.960 ;
        RECT 17.080 99.405 17.310 99.560 ;
        RECT 17.720 99.405 17.950 101.760 ;
        RECT 18.360 100.960 18.590 105.405 ;
        RECT 19.300 104.410 19.700 105.585 ;
        RECT 25.350 104.410 25.700 104.460 ;
        RECT 19.300 104.110 25.700 104.410 ;
        RECT 18.315 99.560 18.775 100.960 ;
        RECT 18.360 99.405 18.590 99.560 ;
        RECT 19.300 99.210 19.700 104.110 ;
        RECT 25.350 104.060 25.700 104.110 ;
        RECT 21.550 103.510 25.700 103.810 ;
        RECT 21.280 103.160 21.510 103.360 ;
        RECT 21.225 101.760 21.685 103.160 ;
        RECT 21.280 99.360 21.510 101.760 ;
        RECT 21.920 100.960 22.150 103.360 ;
        RECT 22.560 103.160 22.790 103.360 ;
        RECT 22.500 101.760 22.960 103.160 ;
        RECT 21.890 99.560 22.350 100.960 ;
        RECT 21.920 99.360 22.150 99.560 ;
        RECT 22.560 99.360 22.790 101.760 ;
        RECT 23.200 100.960 23.430 103.360 ;
        RECT 23.840 103.160 24.070 103.360 ;
        RECT 23.775 101.760 24.235 103.160 ;
        RECT 23.165 99.560 23.625 100.960 ;
        RECT 23.200 99.360 23.430 99.560 ;
        RECT 23.840 99.360 24.070 101.760 ;
        RECT 24.480 100.960 24.710 103.360 ;
        RECT 25.430 102.760 25.700 103.510 ;
        RECT 25.350 102.360 25.700 102.760 ;
        RECT 24.450 99.560 24.810 100.960 ;
        RECT 24.480 99.360 24.710 99.560 ;
        RECT 25.430 99.210 25.700 102.360 ;
        RECT 11.600 98.910 19.700 99.210 ;
        RECT 8.050 97.430 17.300 98.495 ;
        RECT 17.920 98.010 18.150 98.100 ;
        RECT 18.360 98.010 18.590 98.100 ;
        RECT 19.300 98.010 19.700 98.910 ;
        RECT 20.160 98.910 25.700 99.210 ;
        RECT 17.815 97.660 18.175 98.010 ;
        RECT 18.340 97.660 18.700 98.010 ;
        RECT 19.250 97.660 19.750 98.010 ;
        RECT 17.920 97.100 18.150 97.660 ;
        RECT 18.360 97.100 18.590 97.660 ;
        RECT 19.300 97.610 19.700 97.660 ;
        RECT 16.600 96.910 17.050 96.960 ;
        RECT 20.160 96.910 20.560 98.910 ;
        RECT 25.850 98.760 26.200 107.430 ;
        RECT 133.655 107.420 140.840 108.485 ;
        RECT 141.460 108.000 141.690 108.090 ;
        RECT 141.900 108.000 142.130 108.090 ;
        RECT 142.840 108.000 143.240 108.900 ;
        RECT 144.820 108.000 145.050 108.060 ;
        RECT 145.260 108.000 145.490 108.060 ;
        RECT 141.355 107.650 141.715 108.000 ;
        RECT 141.880 107.650 142.240 108.000 ;
        RECT 142.790 107.650 143.290 108.000 ;
        RECT 144.705 107.650 145.065 108.000 ;
        RECT 145.230 107.650 145.590 108.000 ;
        RECT 141.460 107.090 141.690 107.650 ;
        RECT 141.900 107.090 142.130 107.650 ;
        RECT 142.840 107.600 143.240 107.650 ;
        RECT 144.820 107.060 145.050 107.650 ;
        RECT 145.260 107.060 145.490 107.650 ;
        RECT 146.390 106.955 146.690 108.900 ;
        RECT 149.390 108.485 149.740 116.475 ;
        RECT 146.840 107.420 151.990 108.485 ;
        RECT 139.690 106.900 140.090 106.950 ;
        RECT 146.335 106.900 146.745 106.955 ;
        RECT 139.690 106.650 146.745 106.900 ;
        RECT 139.690 106.600 140.090 106.650 ;
        RECT 146.335 106.595 146.745 106.650 ;
        RECT 22.670 98.560 26.200 98.760 ;
        RECT 21.280 98.010 21.510 98.070 ;
        RECT 21.720 98.010 21.950 98.070 ;
        RECT 21.165 97.660 21.525 98.010 ;
        RECT 21.690 97.660 22.050 98.010 ;
        RECT 22.670 97.660 23.200 98.560 ;
        RECT 25.100 98.495 26.200 98.560 ;
        RECT 23.920 98.010 24.150 98.060 ;
        RECT 23.775 97.660 24.150 98.010 ;
        RECT 21.280 97.070 21.510 97.660 ;
        RECT 21.720 97.070 21.950 97.660 ;
        RECT 23.920 97.060 24.150 97.660 ;
        RECT 24.360 98.010 24.590 98.060 ;
        RECT 24.360 97.660 24.740 98.010 ;
        RECT 24.360 97.060 24.590 97.660 ;
        RECT 25.100 97.430 26.335 98.495 ;
        RECT 133.790 98.485 134.140 106.475 ;
        RECT 134.290 105.875 134.640 105.925 ;
        RECT 134.290 105.575 143.240 105.875 ;
        RECT 134.860 103.150 135.090 105.395 ;
        RECT 134.815 101.750 135.275 103.150 ;
        RECT 134.860 99.395 135.090 101.750 ;
        RECT 135.500 100.950 135.730 105.395 ;
        RECT 136.140 103.150 136.370 105.395 ;
        RECT 136.090 101.750 136.550 103.150 ;
        RECT 135.465 99.550 135.925 100.950 ;
        RECT 135.500 99.395 135.730 99.550 ;
        RECT 136.140 99.395 136.370 101.750 ;
        RECT 136.780 100.950 137.010 105.395 ;
        RECT 137.420 103.150 137.650 105.395 ;
        RECT 137.365 101.750 137.825 103.150 ;
        RECT 136.755 99.550 137.215 100.950 ;
        RECT 136.780 99.395 137.010 99.550 ;
        RECT 137.420 99.395 137.650 101.750 ;
        RECT 138.060 100.950 138.290 105.395 ;
        RECT 138.700 103.150 138.930 105.395 ;
        RECT 138.640 101.750 139.100 103.150 ;
        RECT 138.030 99.550 138.490 100.950 ;
        RECT 138.060 99.395 138.290 99.550 ;
        RECT 138.700 99.395 138.930 101.750 ;
        RECT 139.340 100.950 139.570 105.395 ;
        RECT 139.980 103.150 140.210 105.395 ;
        RECT 139.915 101.750 140.375 103.150 ;
        RECT 139.305 99.550 139.765 100.950 ;
        RECT 139.340 99.395 139.570 99.550 ;
        RECT 139.980 99.395 140.210 101.750 ;
        RECT 140.620 100.950 140.850 105.395 ;
        RECT 141.260 103.150 141.490 105.395 ;
        RECT 141.190 101.750 141.650 103.150 ;
        RECT 140.580 99.550 141.040 100.950 ;
        RECT 140.620 99.395 140.850 99.550 ;
        RECT 141.260 99.395 141.490 101.750 ;
        RECT 141.900 100.950 142.130 105.395 ;
        RECT 141.855 99.550 142.315 100.950 ;
        RECT 141.900 99.395 142.130 99.550 ;
        RECT 142.840 99.200 143.240 105.575 ;
        RECT 145.090 103.500 149.240 103.800 ;
        RECT 144.820 103.150 145.050 103.350 ;
        RECT 144.765 101.750 145.225 103.150 ;
        RECT 144.820 99.350 145.050 101.750 ;
        RECT 145.460 100.950 145.690 103.350 ;
        RECT 146.100 103.150 146.330 103.350 ;
        RECT 146.040 101.750 146.500 103.150 ;
        RECT 145.430 99.550 145.890 100.950 ;
        RECT 145.460 99.350 145.690 99.550 ;
        RECT 146.100 99.350 146.330 101.750 ;
        RECT 146.740 100.950 146.970 103.350 ;
        RECT 147.380 103.150 147.610 103.350 ;
        RECT 147.315 101.750 147.775 103.150 ;
        RECT 146.705 99.550 147.165 100.950 ;
        RECT 146.740 99.350 146.970 99.550 ;
        RECT 147.380 99.350 147.610 101.750 ;
        RECT 148.020 100.950 148.250 103.350 ;
        RECT 147.990 99.550 148.350 100.950 ;
        RECT 148.020 99.350 148.250 99.550 ;
        RECT 148.970 99.200 149.240 103.500 ;
        RECT 135.140 98.900 143.240 99.200 ;
        RECT 145.090 98.900 149.240 99.200 ;
        RECT 16.600 96.680 21.760 96.910 ;
        RECT 16.600 96.660 21.735 96.680 ;
        RECT 16.600 96.610 17.050 96.660 ;
        RECT 24.025 96.595 24.475 96.915 ;
        RECT 10.250 88.495 10.600 96.485 ;
        RECT 11.600 95.585 19.700 95.885 ;
        RECT 11.320 93.160 11.550 95.405 ;
        RECT 11.275 91.760 11.735 93.160 ;
        RECT 11.320 89.405 11.550 91.760 ;
        RECT 11.960 90.960 12.190 95.405 ;
        RECT 12.600 93.160 12.830 95.405 ;
        RECT 12.550 91.760 13.010 93.160 ;
        RECT 11.925 89.560 12.385 90.960 ;
        RECT 11.960 89.405 12.190 89.560 ;
        RECT 12.600 89.405 12.830 91.760 ;
        RECT 13.240 90.960 13.470 95.405 ;
        RECT 13.880 93.160 14.110 95.405 ;
        RECT 13.825 91.760 14.285 93.160 ;
        RECT 13.215 89.560 13.675 90.960 ;
        RECT 13.240 89.405 13.470 89.560 ;
        RECT 13.880 89.405 14.110 91.760 ;
        RECT 14.520 90.960 14.750 95.405 ;
        RECT 15.160 93.160 15.390 95.405 ;
        RECT 15.100 91.760 15.560 93.160 ;
        RECT 14.490 89.560 14.950 90.960 ;
        RECT 14.520 89.405 14.750 89.560 ;
        RECT 15.160 89.405 15.390 91.760 ;
        RECT 15.800 90.960 16.030 95.405 ;
        RECT 16.440 93.160 16.670 95.405 ;
        RECT 16.375 91.760 16.835 93.160 ;
        RECT 15.765 89.560 16.225 90.960 ;
        RECT 15.800 89.405 16.030 89.560 ;
        RECT 16.440 89.405 16.670 91.760 ;
        RECT 17.080 90.960 17.310 95.405 ;
        RECT 17.720 93.160 17.950 95.405 ;
        RECT 17.650 91.760 18.110 93.160 ;
        RECT 17.040 89.560 17.500 90.960 ;
        RECT 17.080 89.405 17.310 89.560 ;
        RECT 17.720 89.405 17.950 91.760 ;
        RECT 18.360 90.960 18.590 95.405 ;
        RECT 19.300 94.410 19.700 95.585 ;
        RECT 25.350 94.410 25.700 94.460 ;
        RECT 19.300 94.110 25.700 94.410 ;
        RECT 18.315 89.560 18.775 90.960 ;
        RECT 18.360 89.405 18.590 89.560 ;
        RECT 19.300 89.210 19.700 94.110 ;
        RECT 25.350 94.060 25.700 94.110 ;
        RECT 21.550 93.510 25.700 93.810 ;
        RECT 21.280 93.160 21.510 93.360 ;
        RECT 21.225 91.760 21.685 93.160 ;
        RECT 21.280 89.360 21.510 91.760 ;
        RECT 21.920 90.960 22.150 93.360 ;
        RECT 22.560 93.160 22.790 93.360 ;
        RECT 22.500 91.760 22.960 93.160 ;
        RECT 21.890 89.560 22.350 90.960 ;
        RECT 21.920 89.360 22.150 89.560 ;
        RECT 22.560 89.360 22.790 91.760 ;
        RECT 23.200 90.960 23.430 93.360 ;
        RECT 23.840 93.160 24.070 93.360 ;
        RECT 23.775 91.760 24.235 93.160 ;
        RECT 23.165 89.560 23.625 90.960 ;
        RECT 23.200 89.360 23.430 89.560 ;
        RECT 23.840 89.360 24.070 91.760 ;
        RECT 24.480 90.960 24.710 93.360 ;
        RECT 25.430 92.760 25.700 93.510 ;
        RECT 25.350 92.360 25.700 92.760 ;
        RECT 24.450 89.560 24.810 90.960 ;
        RECT 24.480 89.360 24.710 89.560 ;
        RECT 25.430 89.210 25.700 92.360 ;
        RECT 11.600 88.910 19.700 89.210 ;
        RECT 8.050 87.430 17.300 88.495 ;
        RECT 17.920 88.010 18.150 88.100 ;
        RECT 18.360 88.010 18.590 88.100 ;
        RECT 19.300 88.010 19.700 88.910 ;
        RECT 20.160 88.910 25.700 89.210 ;
        RECT 17.815 87.660 18.175 88.010 ;
        RECT 18.340 87.660 18.700 88.010 ;
        RECT 19.250 87.660 19.750 88.010 ;
        RECT 17.920 87.100 18.150 87.660 ;
        RECT 18.360 87.100 18.590 87.660 ;
        RECT 19.300 87.610 19.700 87.660 ;
        RECT 16.600 86.910 17.050 86.960 ;
        RECT 20.160 86.910 20.560 88.910 ;
        RECT 25.850 88.760 26.200 97.430 ;
        RECT 133.655 97.420 140.840 98.485 ;
        RECT 141.460 98.000 141.690 98.090 ;
        RECT 141.900 98.000 142.130 98.090 ;
        RECT 142.840 98.000 143.240 98.900 ;
        RECT 144.820 98.000 145.050 98.060 ;
        RECT 145.260 98.000 145.490 98.060 ;
        RECT 141.355 97.650 141.715 98.000 ;
        RECT 141.880 97.650 142.240 98.000 ;
        RECT 142.790 97.650 143.290 98.000 ;
        RECT 144.705 97.650 145.065 98.000 ;
        RECT 145.230 97.650 145.590 98.000 ;
        RECT 141.460 97.090 141.690 97.650 ;
        RECT 141.900 97.090 142.130 97.650 ;
        RECT 142.840 97.600 143.240 97.650 ;
        RECT 144.820 97.060 145.050 97.650 ;
        RECT 145.260 97.060 145.490 97.650 ;
        RECT 146.390 96.955 146.690 98.900 ;
        RECT 149.390 98.485 149.740 106.475 ;
        RECT 146.840 97.420 151.990 98.485 ;
        RECT 139.690 96.900 140.090 96.950 ;
        RECT 146.335 96.900 146.745 96.955 ;
        RECT 139.690 96.650 146.745 96.900 ;
        RECT 139.690 96.600 140.090 96.650 ;
        RECT 146.335 96.595 146.745 96.650 ;
        RECT 22.670 88.560 26.200 88.760 ;
        RECT 21.280 88.010 21.510 88.070 ;
        RECT 21.720 88.010 21.950 88.070 ;
        RECT 21.165 87.660 21.525 88.010 ;
        RECT 21.690 87.660 22.050 88.010 ;
        RECT 22.670 87.660 23.200 88.560 ;
        RECT 25.100 88.495 26.200 88.560 ;
        RECT 23.920 88.010 24.150 88.060 ;
        RECT 23.775 87.660 24.150 88.010 ;
        RECT 21.280 87.070 21.510 87.660 ;
        RECT 21.720 87.070 21.950 87.660 ;
        RECT 23.920 87.060 24.150 87.660 ;
        RECT 24.360 88.010 24.590 88.060 ;
        RECT 24.360 87.660 24.740 88.010 ;
        RECT 24.360 87.060 24.590 87.660 ;
        RECT 25.100 87.430 26.335 88.495 ;
        RECT 133.790 88.485 134.140 96.475 ;
        RECT 134.290 95.875 134.640 95.925 ;
        RECT 134.290 95.575 143.240 95.875 ;
        RECT 134.860 93.150 135.090 95.395 ;
        RECT 134.815 91.750 135.275 93.150 ;
        RECT 134.860 89.395 135.090 91.750 ;
        RECT 135.500 90.950 135.730 95.395 ;
        RECT 136.140 93.150 136.370 95.395 ;
        RECT 136.090 91.750 136.550 93.150 ;
        RECT 135.465 89.550 135.925 90.950 ;
        RECT 135.500 89.395 135.730 89.550 ;
        RECT 136.140 89.395 136.370 91.750 ;
        RECT 136.780 90.950 137.010 95.395 ;
        RECT 137.420 93.150 137.650 95.395 ;
        RECT 137.365 91.750 137.825 93.150 ;
        RECT 136.755 89.550 137.215 90.950 ;
        RECT 136.780 89.395 137.010 89.550 ;
        RECT 137.420 89.395 137.650 91.750 ;
        RECT 138.060 90.950 138.290 95.395 ;
        RECT 138.700 93.150 138.930 95.395 ;
        RECT 138.640 91.750 139.100 93.150 ;
        RECT 138.030 89.550 138.490 90.950 ;
        RECT 138.060 89.395 138.290 89.550 ;
        RECT 138.700 89.395 138.930 91.750 ;
        RECT 139.340 90.950 139.570 95.395 ;
        RECT 139.980 93.150 140.210 95.395 ;
        RECT 139.915 91.750 140.375 93.150 ;
        RECT 139.305 89.550 139.765 90.950 ;
        RECT 139.340 89.395 139.570 89.550 ;
        RECT 139.980 89.395 140.210 91.750 ;
        RECT 140.620 90.950 140.850 95.395 ;
        RECT 141.260 93.150 141.490 95.395 ;
        RECT 141.190 91.750 141.650 93.150 ;
        RECT 140.580 89.550 141.040 90.950 ;
        RECT 140.620 89.395 140.850 89.550 ;
        RECT 141.260 89.395 141.490 91.750 ;
        RECT 141.900 90.950 142.130 95.395 ;
        RECT 141.855 89.550 142.315 90.950 ;
        RECT 141.900 89.395 142.130 89.550 ;
        RECT 142.840 89.200 143.240 95.575 ;
        RECT 145.090 93.500 149.240 93.800 ;
        RECT 144.820 93.150 145.050 93.350 ;
        RECT 144.765 91.750 145.225 93.150 ;
        RECT 144.820 89.350 145.050 91.750 ;
        RECT 145.460 90.950 145.690 93.350 ;
        RECT 146.100 93.150 146.330 93.350 ;
        RECT 146.040 91.750 146.500 93.150 ;
        RECT 145.430 89.550 145.890 90.950 ;
        RECT 145.460 89.350 145.690 89.550 ;
        RECT 146.100 89.350 146.330 91.750 ;
        RECT 146.740 90.950 146.970 93.350 ;
        RECT 147.380 93.150 147.610 93.350 ;
        RECT 147.315 91.750 147.775 93.150 ;
        RECT 146.705 89.550 147.165 90.950 ;
        RECT 146.740 89.350 146.970 89.550 ;
        RECT 147.380 89.350 147.610 91.750 ;
        RECT 148.020 90.950 148.250 93.350 ;
        RECT 147.990 89.550 148.350 90.950 ;
        RECT 148.020 89.350 148.250 89.550 ;
        RECT 148.970 89.200 149.240 93.500 ;
        RECT 135.140 88.900 143.240 89.200 ;
        RECT 145.090 88.900 149.240 89.200 ;
        RECT 16.600 86.680 21.760 86.910 ;
        RECT 16.600 86.660 21.735 86.680 ;
        RECT 16.600 86.610 17.050 86.660 ;
        RECT 24.025 86.595 24.475 86.915 ;
        RECT 10.250 78.495 10.600 86.485 ;
        RECT 11.600 85.585 19.700 85.885 ;
        RECT 11.320 83.160 11.550 85.405 ;
        RECT 11.275 81.760 11.735 83.160 ;
        RECT 11.320 79.405 11.550 81.760 ;
        RECT 11.960 80.960 12.190 85.405 ;
        RECT 12.600 83.160 12.830 85.405 ;
        RECT 12.550 81.760 13.010 83.160 ;
        RECT 11.925 79.560 12.385 80.960 ;
        RECT 11.960 79.405 12.190 79.560 ;
        RECT 12.600 79.405 12.830 81.760 ;
        RECT 13.240 80.960 13.470 85.405 ;
        RECT 13.880 83.160 14.110 85.405 ;
        RECT 13.825 81.760 14.285 83.160 ;
        RECT 13.215 79.560 13.675 80.960 ;
        RECT 13.240 79.405 13.470 79.560 ;
        RECT 13.880 79.405 14.110 81.760 ;
        RECT 14.520 80.960 14.750 85.405 ;
        RECT 15.160 83.160 15.390 85.405 ;
        RECT 15.100 81.760 15.560 83.160 ;
        RECT 14.490 79.560 14.950 80.960 ;
        RECT 14.520 79.405 14.750 79.560 ;
        RECT 15.160 79.405 15.390 81.760 ;
        RECT 15.800 80.960 16.030 85.405 ;
        RECT 16.440 83.160 16.670 85.405 ;
        RECT 16.375 81.760 16.835 83.160 ;
        RECT 15.765 79.560 16.225 80.960 ;
        RECT 15.800 79.405 16.030 79.560 ;
        RECT 16.440 79.405 16.670 81.760 ;
        RECT 17.080 80.960 17.310 85.405 ;
        RECT 17.720 83.160 17.950 85.405 ;
        RECT 17.650 81.760 18.110 83.160 ;
        RECT 17.040 79.560 17.500 80.960 ;
        RECT 17.080 79.405 17.310 79.560 ;
        RECT 17.720 79.405 17.950 81.760 ;
        RECT 18.360 80.960 18.590 85.405 ;
        RECT 19.300 84.410 19.700 85.585 ;
        RECT 25.350 84.410 25.700 84.460 ;
        RECT 19.300 84.110 25.700 84.410 ;
        RECT 18.315 79.560 18.775 80.960 ;
        RECT 18.360 79.405 18.590 79.560 ;
        RECT 19.300 79.210 19.700 84.110 ;
        RECT 25.350 84.060 25.700 84.110 ;
        RECT 21.550 83.510 25.700 83.810 ;
        RECT 21.280 83.160 21.510 83.360 ;
        RECT 21.225 81.760 21.685 83.160 ;
        RECT 21.280 79.360 21.510 81.760 ;
        RECT 21.920 80.960 22.150 83.360 ;
        RECT 22.560 83.160 22.790 83.360 ;
        RECT 22.500 81.760 22.960 83.160 ;
        RECT 21.890 79.560 22.350 80.960 ;
        RECT 21.920 79.360 22.150 79.560 ;
        RECT 22.560 79.360 22.790 81.760 ;
        RECT 23.200 80.960 23.430 83.360 ;
        RECT 23.840 83.160 24.070 83.360 ;
        RECT 23.775 81.760 24.235 83.160 ;
        RECT 23.165 79.560 23.625 80.960 ;
        RECT 23.200 79.360 23.430 79.560 ;
        RECT 23.840 79.360 24.070 81.760 ;
        RECT 24.480 80.960 24.710 83.360 ;
        RECT 25.430 82.760 25.700 83.510 ;
        RECT 25.350 82.360 25.700 82.760 ;
        RECT 24.450 79.560 24.810 80.960 ;
        RECT 24.480 79.360 24.710 79.560 ;
        RECT 25.430 79.210 25.700 82.360 ;
        RECT 11.600 78.910 19.700 79.210 ;
        RECT 8.050 77.430 17.300 78.495 ;
        RECT 17.920 78.010 18.150 78.100 ;
        RECT 18.360 78.010 18.590 78.100 ;
        RECT 19.300 78.010 19.700 78.910 ;
        RECT 20.160 78.910 25.700 79.210 ;
        RECT 17.815 77.660 18.175 78.010 ;
        RECT 18.340 77.660 18.700 78.010 ;
        RECT 19.250 77.660 19.750 78.010 ;
        RECT 17.920 77.100 18.150 77.660 ;
        RECT 18.360 77.100 18.590 77.660 ;
        RECT 19.300 77.610 19.700 77.660 ;
        RECT 16.600 76.910 17.050 76.960 ;
        RECT 20.160 76.910 20.560 78.910 ;
        RECT 25.850 78.760 26.200 87.430 ;
        RECT 133.655 87.420 140.840 88.485 ;
        RECT 141.460 88.000 141.690 88.090 ;
        RECT 141.900 88.000 142.130 88.090 ;
        RECT 142.840 88.000 143.240 88.900 ;
        RECT 144.820 88.000 145.050 88.060 ;
        RECT 145.260 88.000 145.490 88.060 ;
        RECT 141.355 87.650 141.715 88.000 ;
        RECT 141.880 87.650 142.240 88.000 ;
        RECT 142.790 87.650 143.290 88.000 ;
        RECT 144.705 87.650 145.065 88.000 ;
        RECT 145.230 87.650 145.590 88.000 ;
        RECT 141.460 87.090 141.690 87.650 ;
        RECT 141.900 87.090 142.130 87.650 ;
        RECT 142.840 87.600 143.240 87.650 ;
        RECT 144.820 87.060 145.050 87.650 ;
        RECT 145.260 87.060 145.490 87.650 ;
        RECT 146.390 86.955 146.690 88.900 ;
        RECT 149.390 88.485 149.740 96.475 ;
        RECT 146.840 87.420 151.990 88.485 ;
        RECT 139.690 86.900 140.090 86.950 ;
        RECT 146.335 86.900 146.745 86.955 ;
        RECT 139.690 86.650 146.745 86.900 ;
        RECT 139.690 86.600 140.090 86.650 ;
        RECT 146.335 86.595 146.745 86.650 ;
        RECT 22.670 78.560 26.200 78.760 ;
        RECT 21.280 78.010 21.510 78.070 ;
        RECT 21.720 78.010 21.950 78.070 ;
        RECT 21.165 77.660 21.525 78.010 ;
        RECT 21.690 77.660 22.050 78.010 ;
        RECT 22.670 77.660 23.200 78.560 ;
        RECT 25.100 78.495 26.200 78.560 ;
        RECT 23.920 78.010 24.150 78.060 ;
        RECT 23.775 77.660 24.150 78.010 ;
        RECT 21.280 77.070 21.510 77.660 ;
        RECT 21.720 77.070 21.950 77.660 ;
        RECT 23.920 77.060 24.150 77.660 ;
        RECT 24.360 78.010 24.590 78.060 ;
        RECT 24.360 77.660 24.740 78.010 ;
        RECT 24.360 77.060 24.590 77.660 ;
        RECT 25.100 77.430 26.335 78.495 ;
        RECT 133.790 78.485 134.140 86.475 ;
        RECT 134.290 85.875 134.640 85.925 ;
        RECT 134.290 85.575 143.240 85.875 ;
        RECT 134.860 83.150 135.090 85.395 ;
        RECT 134.815 81.750 135.275 83.150 ;
        RECT 134.860 79.395 135.090 81.750 ;
        RECT 135.500 80.950 135.730 85.395 ;
        RECT 136.140 83.150 136.370 85.395 ;
        RECT 136.090 81.750 136.550 83.150 ;
        RECT 135.465 79.550 135.925 80.950 ;
        RECT 135.500 79.395 135.730 79.550 ;
        RECT 136.140 79.395 136.370 81.750 ;
        RECT 136.780 80.950 137.010 85.395 ;
        RECT 137.420 83.150 137.650 85.395 ;
        RECT 137.365 81.750 137.825 83.150 ;
        RECT 136.755 79.550 137.215 80.950 ;
        RECT 136.780 79.395 137.010 79.550 ;
        RECT 137.420 79.395 137.650 81.750 ;
        RECT 138.060 80.950 138.290 85.395 ;
        RECT 138.700 83.150 138.930 85.395 ;
        RECT 138.640 81.750 139.100 83.150 ;
        RECT 138.030 79.550 138.490 80.950 ;
        RECT 138.060 79.395 138.290 79.550 ;
        RECT 138.700 79.395 138.930 81.750 ;
        RECT 139.340 80.950 139.570 85.395 ;
        RECT 139.980 83.150 140.210 85.395 ;
        RECT 139.915 81.750 140.375 83.150 ;
        RECT 139.305 79.550 139.765 80.950 ;
        RECT 139.340 79.395 139.570 79.550 ;
        RECT 139.980 79.395 140.210 81.750 ;
        RECT 140.620 80.950 140.850 85.395 ;
        RECT 141.260 83.150 141.490 85.395 ;
        RECT 141.190 81.750 141.650 83.150 ;
        RECT 140.580 79.550 141.040 80.950 ;
        RECT 140.620 79.395 140.850 79.550 ;
        RECT 141.260 79.395 141.490 81.750 ;
        RECT 141.900 80.950 142.130 85.395 ;
        RECT 141.855 79.550 142.315 80.950 ;
        RECT 141.900 79.395 142.130 79.550 ;
        RECT 142.840 79.200 143.240 85.575 ;
        RECT 145.090 83.500 149.240 83.800 ;
        RECT 144.820 83.150 145.050 83.350 ;
        RECT 144.765 81.750 145.225 83.150 ;
        RECT 144.820 79.350 145.050 81.750 ;
        RECT 145.460 80.950 145.690 83.350 ;
        RECT 146.100 83.150 146.330 83.350 ;
        RECT 146.040 81.750 146.500 83.150 ;
        RECT 145.430 79.550 145.890 80.950 ;
        RECT 145.460 79.350 145.690 79.550 ;
        RECT 146.100 79.350 146.330 81.750 ;
        RECT 146.740 80.950 146.970 83.350 ;
        RECT 147.380 83.150 147.610 83.350 ;
        RECT 147.315 81.750 147.775 83.150 ;
        RECT 146.705 79.550 147.165 80.950 ;
        RECT 146.740 79.350 146.970 79.550 ;
        RECT 147.380 79.350 147.610 81.750 ;
        RECT 148.020 80.950 148.250 83.350 ;
        RECT 147.990 79.550 148.350 80.950 ;
        RECT 148.020 79.350 148.250 79.550 ;
        RECT 148.970 79.200 149.240 83.500 ;
        RECT 135.140 78.900 143.240 79.200 ;
        RECT 145.090 78.900 149.240 79.200 ;
        RECT 16.600 76.680 21.760 76.910 ;
        RECT 16.600 76.660 21.735 76.680 ;
        RECT 16.600 76.610 17.050 76.660 ;
        RECT 24.025 76.595 24.475 76.915 ;
        RECT 10.250 68.495 10.600 76.485 ;
        RECT 11.600 75.585 19.700 75.885 ;
        RECT 11.320 73.160 11.550 75.405 ;
        RECT 11.275 71.760 11.735 73.160 ;
        RECT 11.320 69.405 11.550 71.760 ;
        RECT 11.960 70.960 12.190 75.405 ;
        RECT 12.600 73.160 12.830 75.405 ;
        RECT 12.550 71.760 13.010 73.160 ;
        RECT 11.925 69.560 12.385 70.960 ;
        RECT 11.960 69.405 12.190 69.560 ;
        RECT 12.600 69.405 12.830 71.760 ;
        RECT 13.240 70.960 13.470 75.405 ;
        RECT 13.880 73.160 14.110 75.405 ;
        RECT 13.825 71.760 14.285 73.160 ;
        RECT 13.215 69.560 13.675 70.960 ;
        RECT 13.240 69.405 13.470 69.560 ;
        RECT 13.880 69.405 14.110 71.760 ;
        RECT 14.520 70.960 14.750 75.405 ;
        RECT 15.160 73.160 15.390 75.405 ;
        RECT 15.100 71.760 15.560 73.160 ;
        RECT 14.490 69.560 14.950 70.960 ;
        RECT 14.520 69.405 14.750 69.560 ;
        RECT 15.160 69.405 15.390 71.760 ;
        RECT 15.800 70.960 16.030 75.405 ;
        RECT 16.440 73.160 16.670 75.405 ;
        RECT 16.375 71.760 16.835 73.160 ;
        RECT 15.765 69.560 16.225 70.960 ;
        RECT 15.800 69.405 16.030 69.560 ;
        RECT 16.440 69.405 16.670 71.760 ;
        RECT 17.080 70.960 17.310 75.405 ;
        RECT 17.720 73.160 17.950 75.405 ;
        RECT 17.650 71.760 18.110 73.160 ;
        RECT 17.040 69.560 17.500 70.960 ;
        RECT 17.080 69.405 17.310 69.560 ;
        RECT 17.720 69.405 17.950 71.760 ;
        RECT 18.360 70.960 18.590 75.405 ;
        RECT 19.300 74.410 19.700 75.585 ;
        RECT 25.350 74.410 25.700 74.460 ;
        RECT 19.300 74.110 25.700 74.410 ;
        RECT 18.315 69.560 18.775 70.960 ;
        RECT 18.360 69.405 18.590 69.560 ;
        RECT 19.300 69.210 19.700 74.110 ;
        RECT 25.350 74.060 25.700 74.110 ;
        RECT 21.550 73.510 25.700 73.810 ;
        RECT 21.280 73.160 21.510 73.360 ;
        RECT 21.225 71.760 21.685 73.160 ;
        RECT 21.280 69.360 21.510 71.760 ;
        RECT 21.920 70.960 22.150 73.360 ;
        RECT 22.560 73.160 22.790 73.360 ;
        RECT 22.500 71.760 22.960 73.160 ;
        RECT 21.890 69.560 22.350 70.960 ;
        RECT 21.920 69.360 22.150 69.560 ;
        RECT 22.560 69.360 22.790 71.760 ;
        RECT 23.200 70.960 23.430 73.360 ;
        RECT 23.840 73.160 24.070 73.360 ;
        RECT 23.775 71.760 24.235 73.160 ;
        RECT 23.165 69.560 23.625 70.960 ;
        RECT 23.200 69.360 23.430 69.560 ;
        RECT 23.840 69.360 24.070 71.760 ;
        RECT 24.480 70.960 24.710 73.360 ;
        RECT 25.430 72.760 25.700 73.510 ;
        RECT 25.350 72.360 25.700 72.760 ;
        RECT 24.450 69.560 24.810 70.960 ;
        RECT 24.480 69.360 24.710 69.560 ;
        RECT 25.430 69.210 25.700 72.360 ;
        RECT 11.600 68.910 19.700 69.210 ;
        RECT 8.050 67.430 17.300 68.495 ;
        RECT 17.920 68.010 18.150 68.100 ;
        RECT 18.360 68.010 18.590 68.100 ;
        RECT 19.300 68.010 19.700 68.910 ;
        RECT 20.160 68.910 25.700 69.210 ;
        RECT 17.815 67.660 18.175 68.010 ;
        RECT 18.340 67.660 18.700 68.010 ;
        RECT 19.250 67.660 19.750 68.010 ;
        RECT 17.920 67.100 18.150 67.660 ;
        RECT 18.360 67.100 18.590 67.660 ;
        RECT 19.300 67.610 19.700 67.660 ;
        RECT 16.600 66.910 17.050 66.960 ;
        RECT 20.160 66.910 20.560 68.910 ;
        RECT 25.850 68.760 26.200 77.430 ;
        RECT 133.655 77.420 140.840 78.485 ;
        RECT 141.460 78.000 141.690 78.090 ;
        RECT 141.900 78.000 142.130 78.090 ;
        RECT 142.840 78.000 143.240 78.900 ;
        RECT 144.820 78.000 145.050 78.060 ;
        RECT 145.260 78.000 145.490 78.060 ;
        RECT 141.355 77.650 141.715 78.000 ;
        RECT 141.880 77.650 142.240 78.000 ;
        RECT 142.790 77.650 143.290 78.000 ;
        RECT 144.705 77.650 145.065 78.000 ;
        RECT 145.230 77.650 145.590 78.000 ;
        RECT 141.460 77.090 141.690 77.650 ;
        RECT 141.900 77.090 142.130 77.650 ;
        RECT 142.840 77.600 143.240 77.650 ;
        RECT 144.820 77.060 145.050 77.650 ;
        RECT 145.260 77.060 145.490 77.650 ;
        RECT 146.390 76.955 146.690 78.900 ;
        RECT 149.390 78.485 149.740 86.475 ;
        RECT 146.840 77.420 151.990 78.485 ;
        RECT 139.690 76.900 140.090 76.950 ;
        RECT 146.335 76.900 146.745 76.955 ;
        RECT 139.690 76.650 146.745 76.900 ;
        RECT 139.690 76.600 140.090 76.650 ;
        RECT 146.335 76.595 146.745 76.650 ;
        RECT 22.670 68.560 26.200 68.760 ;
        RECT 21.280 68.010 21.510 68.070 ;
        RECT 21.720 68.010 21.950 68.070 ;
        RECT 21.165 67.660 21.525 68.010 ;
        RECT 21.690 67.660 22.050 68.010 ;
        RECT 22.670 67.660 23.200 68.560 ;
        RECT 25.100 68.495 26.200 68.560 ;
        RECT 23.920 68.010 24.150 68.060 ;
        RECT 23.775 67.660 24.150 68.010 ;
        RECT 21.280 67.070 21.510 67.660 ;
        RECT 21.720 67.070 21.950 67.660 ;
        RECT 23.920 67.060 24.150 67.660 ;
        RECT 24.360 68.010 24.590 68.060 ;
        RECT 24.360 67.660 24.740 68.010 ;
        RECT 24.360 67.060 24.590 67.660 ;
        RECT 25.100 67.430 26.335 68.495 ;
        RECT 133.790 68.485 134.140 76.475 ;
        RECT 134.290 75.875 134.640 75.925 ;
        RECT 134.290 75.575 143.240 75.875 ;
        RECT 134.860 73.150 135.090 75.395 ;
        RECT 134.815 71.750 135.275 73.150 ;
        RECT 134.860 69.395 135.090 71.750 ;
        RECT 135.500 70.950 135.730 75.395 ;
        RECT 136.140 73.150 136.370 75.395 ;
        RECT 136.090 71.750 136.550 73.150 ;
        RECT 135.465 69.550 135.925 70.950 ;
        RECT 135.500 69.395 135.730 69.550 ;
        RECT 136.140 69.395 136.370 71.750 ;
        RECT 136.780 70.950 137.010 75.395 ;
        RECT 137.420 73.150 137.650 75.395 ;
        RECT 137.365 71.750 137.825 73.150 ;
        RECT 136.755 69.550 137.215 70.950 ;
        RECT 136.780 69.395 137.010 69.550 ;
        RECT 137.420 69.395 137.650 71.750 ;
        RECT 138.060 70.950 138.290 75.395 ;
        RECT 138.700 73.150 138.930 75.395 ;
        RECT 138.640 71.750 139.100 73.150 ;
        RECT 138.030 69.550 138.490 70.950 ;
        RECT 138.060 69.395 138.290 69.550 ;
        RECT 138.700 69.395 138.930 71.750 ;
        RECT 139.340 70.950 139.570 75.395 ;
        RECT 139.980 73.150 140.210 75.395 ;
        RECT 139.915 71.750 140.375 73.150 ;
        RECT 139.305 69.550 139.765 70.950 ;
        RECT 139.340 69.395 139.570 69.550 ;
        RECT 139.980 69.395 140.210 71.750 ;
        RECT 140.620 70.950 140.850 75.395 ;
        RECT 141.260 73.150 141.490 75.395 ;
        RECT 141.190 71.750 141.650 73.150 ;
        RECT 140.580 69.550 141.040 70.950 ;
        RECT 140.620 69.395 140.850 69.550 ;
        RECT 141.260 69.395 141.490 71.750 ;
        RECT 141.900 70.950 142.130 75.395 ;
        RECT 141.855 69.550 142.315 70.950 ;
        RECT 141.900 69.395 142.130 69.550 ;
        RECT 142.840 69.200 143.240 75.575 ;
        RECT 145.090 73.500 149.240 73.800 ;
        RECT 144.820 73.150 145.050 73.350 ;
        RECT 144.765 71.750 145.225 73.150 ;
        RECT 144.820 69.350 145.050 71.750 ;
        RECT 145.460 70.950 145.690 73.350 ;
        RECT 146.100 73.150 146.330 73.350 ;
        RECT 146.040 71.750 146.500 73.150 ;
        RECT 145.430 69.550 145.890 70.950 ;
        RECT 145.460 69.350 145.690 69.550 ;
        RECT 146.100 69.350 146.330 71.750 ;
        RECT 146.740 70.950 146.970 73.350 ;
        RECT 147.380 73.150 147.610 73.350 ;
        RECT 147.315 71.750 147.775 73.150 ;
        RECT 146.705 69.550 147.165 70.950 ;
        RECT 146.740 69.350 146.970 69.550 ;
        RECT 147.380 69.350 147.610 71.750 ;
        RECT 148.020 70.950 148.250 73.350 ;
        RECT 147.990 69.550 148.350 70.950 ;
        RECT 148.020 69.350 148.250 69.550 ;
        RECT 148.970 69.200 149.240 73.500 ;
        RECT 135.140 68.900 143.240 69.200 ;
        RECT 145.090 68.900 149.240 69.200 ;
        RECT 16.600 66.680 21.760 66.910 ;
        RECT 16.600 66.660 21.735 66.680 ;
        RECT 16.600 66.610 17.050 66.660 ;
        RECT 24.025 66.595 24.475 66.915 ;
        RECT 10.250 58.495 10.600 66.485 ;
        RECT 11.600 65.585 19.700 65.885 ;
        RECT 11.320 63.160 11.550 65.405 ;
        RECT 11.275 61.760 11.735 63.160 ;
        RECT 11.320 59.405 11.550 61.760 ;
        RECT 11.960 60.960 12.190 65.405 ;
        RECT 12.600 63.160 12.830 65.405 ;
        RECT 12.550 61.760 13.010 63.160 ;
        RECT 11.925 59.560 12.385 60.960 ;
        RECT 11.960 59.405 12.190 59.560 ;
        RECT 12.600 59.405 12.830 61.760 ;
        RECT 13.240 60.960 13.470 65.405 ;
        RECT 13.880 63.160 14.110 65.405 ;
        RECT 13.825 61.760 14.285 63.160 ;
        RECT 13.215 59.560 13.675 60.960 ;
        RECT 13.240 59.405 13.470 59.560 ;
        RECT 13.880 59.405 14.110 61.760 ;
        RECT 14.520 60.960 14.750 65.405 ;
        RECT 15.160 63.160 15.390 65.405 ;
        RECT 15.100 61.760 15.560 63.160 ;
        RECT 14.490 59.560 14.950 60.960 ;
        RECT 14.520 59.405 14.750 59.560 ;
        RECT 15.160 59.405 15.390 61.760 ;
        RECT 15.800 60.960 16.030 65.405 ;
        RECT 16.440 63.160 16.670 65.405 ;
        RECT 16.375 61.760 16.835 63.160 ;
        RECT 15.765 59.560 16.225 60.960 ;
        RECT 15.800 59.405 16.030 59.560 ;
        RECT 16.440 59.405 16.670 61.760 ;
        RECT 17.080 60.960 17.310 65.405 ;
        RECT 17.720 63.160 17.950 65.405 ;
        RECT 17.650 61.760 18.110 63.160 ;
        RECT 17.040 59.560 17.500 60.960 ;
        RECT 17.080 59.405 17.310 59.560 ;
        RECT 17.720 59.405 17.950 61.760 ;
        RECT 18.360 60.960 18.590 65.405 ;
        RECT 19.300 64.410 19.700 65.585 ;
        RECT 25.350 64.410 25.700 64.460 ;
        RECT 19.300 64.110 25.700 64.410 ;
        RECT 18.315 59.560 18.775 60.960 ;
        RECT 18.360 59.405 18.590 59.560 ;
        RECT 19.300 59.210 19.700 64.110 ;
        RECT 25.350 64.060 25.700 64.110 ;
        RECT 21.550 63.510 25.700 63.810 ;
        RECT 21.280 63.160 21.510 63.360 ;
        RECT 21.225 61.760 21.685 63.160 ;
        RECT 21.280 59.360 21.510 61.760 ;
        RECT 21.920 60.960 22.150 63.360 ;
        RECT 22.560 63.160 22.790 63.360 ;
        RECT 22.500 61.760 22.960 63.160 ;
        RECT 21.890 59.560 22.350 60.960 ;
        RECT 21.920 59.360 22.150 59.560 ;
        RECT 22.560 59.360 22.790 61.760 ;
        RECT 23.200 60.960 23.430 63.360 ;
        RECT 23.840 63.160 24.070 63.360 ;
        RECT 23.775 61.760 24.235 63.160 ;
        RECT 23.165 59.560 23.625 60.960 ;
        RECT 23.200 59.360 23.430 59.560 ;
        RECT 23.840 59.360 24.070 61.760 ;
        RECT 24.480 60.960 24.710 63.360 ;
        RECT 25.430 62.760 25.700 63.510 ;
        RECT 25.350 62.360 25.700 62.760 ;
        RECT 24.450 59.560 24.810 60.960 ;
        RECT 24.480 59.360 24.710 59.560 ;
        RECT 25.430 59.210 25.700 62.360 ;
        RECT 11.600 58.910 19.700 59.210 ;
        RECT 8.050 57.430 17.300 58.495 ;
        RECT 17.920 58.010 18.150 58.100 ;
        RECT 18.360 58.010 18.590 58.100 ;
        RECT 19.300 58.010 19.700 58.910 ;
        RECT 20.160 58.910 25.700 59.210 ;
        RECT 17.815 57.660 18.175 58.010 ;
        RECT 18.340 57.660 18.700 58.010 ;
        RECT 19.250 57.660 19.750 58.010 ;
        RECT 17.920 57.100 18.150 57.660 ;
        RECT 18.360 57.100 18.590 57.660 ;
        RECT 19.300 57.610 19.700 57.660 ;
        RECT 16.600 56.910 17.050 56.960 ;
        RECT 20.160 56.910 20.560 58.910 ;
        RECT 25.850 58.760 26.200 67.430 ;
        RECT 133.655 67.420 140.840 68.485 ;
        RECT 141.460 68.000 141.690 68.090 ;
        RECT 141.900 68.000 142.130 68.090 ;
        RECT 142.840 68.000 143.240 68.900 ;
        RECT 144.820 68.000 145.050 68.060 ;
        RECT 145.260 68.000 145.490 68.060 ;
        RECT 141.355 67.650 141.715 68.000 ;
        RECT 141.880 67.650 142.240 68.000 ;
        RECT 142.790 67.650 143.290 68.000 ;
        RECT 144.705 67.650 145.065 68.000 ;
        RECT 145.230 67.650 145.590 68.000 ;
        RECT 141.460 67.090 141.690 67.650 ;
        RECT 141.900 67.090 142.130 67.650 ;
        RECT 142.840 67.600 143.240 67.650 ;
        RECT 144.820 67.060 145.050 67.650 ;
        RECT 145.260 67.060 145.490 67.650 ;
        RECT 146.390 66.955 146.690 68.900 ;
        RECT 149.390 68.485 149.740 76.475 ;
        RECT 146.840 67.420 151.990 68.485 ;
        RECT 139.690 66.900 140.090 66.950 ;
        RECT 146.335 66.900 146.745 66.955 ;
        RECT 139.690 66.650 146.745 66.900 ;
        RECT 139.690 66.600 140.090 66.650 ;
        RECT 146.335 66.595 146.745 66.650 ;
        RECT 22.670 58.560 26.200 58.760 ;
        RECT 21.280 58.010 21.510 58.070 ;
        RECT 21.720 58.010 21.950 58.070 ;
        RECT 21.165 57.660 21.525 58.010 ;
        RECT 21.690 57.660 22.050 58.010 ;
        RECT 22.670 57.660 23.200 58.560 ;
        RECT 25.100 58.495 26.200 58.560 ;
        RECT 23.920 58.010 24.150 58.060 ;
        RECT 23.775 57.660 24.150 58.010 ;
        RECT 21.280 57.070 21.510 57.660 ;
        RECT 21.720 57.070 21.950 57.660 ;
        RECT 23.920 57.060 24.150 57.660 ;
        RECT 24.360 58.010 24.590 58.060 ;
        RECT 24.360 57.660 24.740 58.010 ;
        RECT 24.360 57.060 24.590 57.660 ;
        RECT 25.100 57.430 26.335 58.495 ;
        RECT 133.790 58.485 134.140 66.475 ;
        RECT 134.290 65.875 134.640 65.925 ;
        RECT 134.290 65.575 143.240 65.875 ;
        RECT 134.860 63.150 135.090 65.395 ;
        RECT 134.815 61.750 135.275 63.150 ;
        RECT 134.860 59.395 135.090 61.750 ;
        RECT 135.500 60.950 135.730 65.395 ;
        RECT 136.140 63.150 136.370 65.395 ;
        RECT 136.090 61.750 136.550 63.150 ;
        RECT 135.465 59.550 135.925 60.950 ;
        RECT 135.500 59.395 135.730 59.550 ;
        RECT 136.140 59.395 136.370 61.750 ;
        RECT 136.780 60.950 137.010 65.395 ;
        RECT 137.420 63.150 137.650 65.395 ;
        RECT 137.365 61.750 137.825 63.150 ;
        RECT 136.755 59.550 137.215 60.950 ;
        RECT 136.780 59.395 137.010 59.550 ;
        RECT 137.420 59.395 137.650 61.750 ;
        RECT 138.060 60.950 138.290 65.395 ;
        RECT 138.700 63.150 138.930 65.395 ;
        RECT 138.640 61.750 139.100 63.150 ;
        RECT 138.030 59.550 138.490 60.950 ;
        RECT 138.060 59.395 138.290 59.550 ;
        RECT 138.700 59.395 138.930 61.750 ;
        RECT 139.340 60.950 139.570 65.395 ;
        RECT 139.980 63.150 140.210 65.395 ;
        RECT 139.915 61.750 140.375 63.150 ;
        RECT 139.305 59.550 139.765 60.950 ;
        RECT 139.340 59.395 139.570 59.550 ;
        RECT 139.980 59.395 140.210 61.750 ;
        RECT 140.620 60.950 140.850 65.395 ;
        RECT 141.260 63.150 141.490 65.395 ;
        RECT 141.190 61.750 141.650 63.150 ;
        RECT 140.580 59.550 141.040 60.950 ;
        RECT 140.620 59.395 140.850 59.550 ;
        RECT 141.260 59.395 141.490 61.750 ;
        RECT 141.900 60.950 142.130 65.395 ;
        RECT 141.855 59.550 142.315 60.950 ;
        RECT 141.900 59.395 142.130 59.550 ;
        RECT 142.840 59.200 143.240 65.575 ;
        RECT 145.090 63.500 149.240 63.800 ;
        RECT 144.820 63.150 145.050 63.350 ;
        RECT 144.765 61.750 145.225 63.150 ;
        RECT 144.820 59.350 145.050 61.750 ;
        RECT 145.460 60.950 145.690 63.350 ;
        RECT 146.100 63.150 146.330 63.350 ;
        RECT 146.040 61.750 146.500 63.150 ;
        RECT 145.430 59.550 145.890 60.950 ;
        RECT 145.460 59.350 145.690 59.550 ;
        RECT 146.100 59.350 146.330 61.750 ;
        RECT 146.740 60.950 146.970 63.350 ;
        RECT 147.380 63.150 147.610 63.350 ;
        RECT 147.315 61.750 147.775 63.150 ;
        RECT 146.705 59.550 147.165 60.950 ;
        RECT 146.740 59.350 146.970 59.550 ;
        RECT 147.380 59.350 147.610 61.750 ;
        RECT 148.020 60.950 148.250 63.350 ;
        RECT 147.990 59.550 148.350 60.950 ;
        RECT 148.020 59.350 148.250 59.550 ;
        RECT 148.970 59.200 149.240 63.500 ;
        RECT 135.140 58.900 143.240 59.200 ;
        RECT 145.090 58.900 149.240 59.200 ;
        RECT 16.600 56.680 21.760 56.910 ;
        RECT 16.600 56.660 21.735 56.680 ;
        RECT 16.600 56.610 17.050 56.660 ;
        RECT 24.025 56.595 24.475 56.915 ;
        RECT 10.250 48.495 10.600 56.485 ;
        RECT 11.600 55.585 19.700 55.885 ;
        RECT 11.320 53.160 11.550 55.405 ;
        RECT 11.275 51.760 11.735 53.160 ;
        RECT 11.320 49.405 11.550 51.760 ;
        RECT 11.960 50.960 12.190 55.405 ;
        RECT 12.600 53.160 12.830 55.405 ;
        RECT 12.550 51.760 13.010 53.160 ;
        RECT 11.925 49.560 12.385 50.960 ;
        RECT 11.960 49.405 12.190 49.560 ;
        RECT 12.600 49.405 12.830 51.760 ;
        RECT 13.240 50.960 13.470 55.405 ;
        RECT 13.880 53.160 14.110 55.405 ;
        RECT 13.825 51.760 14.285 53.160 ;
        RECT 13.215 49.560 13.675 50.960 ;
        RECT 13.240 49.405 13.470 49.560 ;
        RECT 13.880 49.405 14.110 51.760 ;
        RECT 14.520 50.960 14.750 55.405 ;
        RECT 15.160 53.160 15.390 55.405 ;
        RECT 15.100 51.760 15.560 53.160 ;
        RECT 14.490 49.560 14.950 50.960 ;
        RECT 14.520 49.405 14.750 49.560 ;
        RECT 15.160 49.405 15.390 51.760 ;
        RECT 15.800 50.960 16.030 55.405 ;
        RECT 16.440 53.160 16.670 55.405 ;
        RECT 16.375 51.760 16.835 53.160 ;
        RECT 15.765 49.560 16.225 50.960 ;
        RECT 15.800 49.405 16.030 49.560 ;
        RECT 16.440 49.405 16.670 51.760 ;
        RECT 17.080 50.960 17.310 55.405 ;
        RECT 17.720 53.160 17.950 55.405 ;
        RECT 17.650 51.760 18.110 53.160 ;
        RECT 17.040 49.560 17.500 50.960 ;
        RECT 17.080 49.405 17.310 49.560 ;
        RECT 17.720 49.405 17.950 51.760 ;
        RECT 18.360 50.960 18.590 55.405 ;
        RECT 19.300 54.410 19.700 55.585 ;
        RECT 25.350 54.410 25.700 54.460 ;
        RECT 19.300 54.110 25.700 54.410 ;
        RECT 18.315 49.560 18.775 50.960 ;
        RECT 18.360 49.405 18.590 49.560 ;
        RECT 19.300 49.210 19.700 54.110 ;
        RECT 25.350 54.060 25.700 54.110 ;
        RECT 21.550 53.510 25.700 53.810 ;
        RECT 21.280 53.160 21.510 53.360 ;
        RECT 21.225 51.760 21.685 53.160 ;
        RECT 21.280 49.360 21.510 51.760 ;
        RECT 21.920 50.960 22.150 53.360 ;
        RECT 22.560 53.160 22.790 53.360 ;
        RECT 22.500 51.760 22.960 53.160 ;
        RECT 21.890 49.560 22.350 50.960 ;
        RECT 21.920 49.360 22.150 49.560 ;
        RECT 22.560 49.360 22.790 51.760 ;
        RECT 23.200 50.960 23.430 53.360 ;
        RECT 23.840 53.160 24.070 53.360 ;
        RECT 23.775 51.760 24.235 53.160 ;
        RECT 23.165 49.560 23.625 50.960 ;
        RECT 23.200 49.360 23.430 49.560 ;
        RECT 23.840 49.360 24.070 51.760 ;
        RECT 24.480 50.960 24.710 53.360 ;
        RECT 25.430 52.760 25.700 53.510 ;
        RECT 25.350 52.360 25.700 52.760 ;
        RECT 24.450 49.560 24.810 50.960 ;
        RECT 24.480 49.360 24.710 49.560 ;
        RECT 25.430 49.210 25.700 52.360 ;
        RECT 11.600 48.910 19.700 49.210 ;
        RECT 8.050 47.430 17.300 48.495 ;
        RECT 17.920 48.010 18.150 48.100 ;
        RECT 18.360 48.010 18.590 48.100 ;
        RECT 19.300 48.010 19.700 48.910 ;
        RECT 20.160 48.910 25.700 49.210 ;
        RECT 17.815 47.660 18.175 48.010 ;
        RECT 18.340 47.660 18.700 48.010 ;
        RECT 19.250 47.660 19.750 48.010 ;
        RECT 17.920 47.100 18.150 47.660 ;
        RECT 18.360 47.100 18.590 47.660 ;
        RECT 19.300 47.610 19.700 47.660 ;
        RECT 16.600 46.910 17.050 46.960 ;
        RECT 20.160 46.910 20.560 48.910 ;
        RECT 25.850 48.760 26.200 57.430 ;
        RECT 133.655 57.420 140.840 58.485 ;
        RECT 141.460 58.000 141.690 58.090 ;
        RECT 141.900 58.000 142.130 58.090 ;
        RECT 142.840 58.000 143.240 58.900 ;
        RECT 144.820 58.000 145.050 58.060 ;
        RECT 145.260 58.000 145.490 58.060 ;
        RECT 141.355 57.650 141.715 58.000 ;
        RECT 141.880 57.650 142.240 58.000 ;
        RECT 142.790 57.650 143.290 58.000 ;
        RECT 144.705 57.650 145.065 58.000 ;
        RECT 145.230 57.650 145.590 58.000 ;
        RECT 141.460 57.090 141.690 57.650 ;
        RECT 141.900 57.090 142.130 57.650 ;
        RECT 142.840 57.600 143.240 57.650 ;
        RECT 144.820 57.060 145.050 57.650 ;
        RECT 145.260 57.060 145.490 57.650 ;
        RECT 146.390 56.955 146.690 58.900 ;
        RECT 149.390 58.485 149.740 66.475 ;
        RECT 146.840 57.420 151.990 58.485 ;
        RECT 139.690 56.900 140.090 56.950 ;
        RECT 146.335 56.900 146.745 56.955 ;
        RECT 139.690 56.650 146.745 56.900 ;
        RECT 139.690 56.600 140.090 56.650 ;
        RECT 146.335 56.595 146.745 56.650 ;
        RECT 22.670 48.560 26.200 48.760 ;
        RECT 21.280 48.010 21.510 48.070 ;
        RECT 21.720 48.010 21.950 48.070 ;
        RECT 21.165 47.660 21.525 48.010 ;
        RECT 21.690 47.660 22.050 48.010 ;
        RECT 22.670 47.660 23.200 48.560 ;
        RECT 25.100 48.495 26.200 48.560 ;
        RECT 23.920 48.010 24.150 48.060 ;
        RECT 23.775 47.660 24.150 48.010 ;
        RECT 21.280 47.070 21.510 47.660 ;
        RECT 21.720 47.070 21.950 47.660 ;
        RECT 23.920 47.060 24.150 47.660 ;
        RECT 24.360 48.010 24.590 48.060 ;
        RECT 24.360 47.660 24.740 48.010 ;
        RECT 24.360 47.060 24.590 47.660 ;
        RECT 25.100 47.430 26.335 48.495 ;
        RECT 133.790 48.485 134.140 56.475 ;
        RECT 134.290 55.875 134.640 55.925 ;
        RECT 134.290 55.575 143.240 55.875 ;
        RECT 134.860 53.150 135.090 55.395 ;
        RECT 134.815 51.750 135.275 53.150 ;
        RECT 134.860 49.395 135.090 51.750 ;
        RECT 135.500 50.950 135.730 55.395 ;
        RECT 136.140 53.150 136.370 55.395 ;
        RECT 136.090 51.750 136.550 53.150 ;
        RECT 135.465 49.550 135.925 50.950 ;
        RECT 135.500 49.395 135.730 49.550 ;
        RECT 136.140 49.395 136.370 51.750 ;
        RECT 136.780 50.950 137.010 55.395 ;
        RECT 137.420 53.150 137.650 55.395 ;
        RECT 137.365 51.750 137.825 53.150 ;
        RECT 136.755 49.550 137.215 50.950 ;
        RECT 136.780 49.395 137.010 49.550 ;
        RECT 137.420 49.395 137.650 51.750 ;
        RECT 138.060 50.950 138.290 55.395 ;
        RECT 138.700 53.150 138.930 55.395 ;
        RECT 138.640 51.750 139.100 53.150 ;
        RECT 138.030 49.550 138.490 50.950 ;
        RECT 138.060 49.395 138.290 49.550 ;
        RECT 138.700 49.395 138.930 51.750 ;
        RECT 139.340 50.950 139.570 55.395 ;
        RECT 139.980 53.150 140.210 55.395 ;
        RECT 139.915 51.750 140.375 53.150 ;
        RECT 139.305 49.550 139.765 50.950 ;
        RECT 139.340 49.395 139.570 49.550 ;
        RECT 139.980 49.395 140.210 51.750 ;
        RECT 140.620 50.950 140.850 55.395 ;
        RECT 141.260 53.150 141.490 55.395 ;
        RECT 141.190 51.750 141.650 53.150 ;
        RECT 140.580 49.550 141.040 50.950 ;
        RECT 140.620 49.395 140.850 49.550 ;
        RECT 141.260 49.395 141.490 51.750 ;
        RECT 141.900 50.950 142.130 55.395 ;
        RECT 141.855 49.550 142.315 50.950 ;
        RECT 141.900 49.395 142.130 49.550 ;
        RECT 142.840 49.200 143.240 55.575 ;
        RECT 145.090 53.500 149.240 53.800 ;
        RECT 144.820 53.150 145.050 53.350 ;
        RECT 144.765 51.750 145.225 53.150 ;
        RECT 144.820 49.350 145.050 51.750 ;
        RECT 145.460 50.950 145.690 53.350 ;
        RECT 146.100 53.150 146.330 53.350 ;
        RECT 146.040 51.750 146.500 53.150 ;
        RECT 145.430 49.550 145.890 50.950 ;
        RECT 145.460 49.350 145.690 49.550 ;
        RECT 146.100 49.350 146.330 51.750 ;
        RECT 146.740 50.950 146.970 53.350 ;
        RECT 147.380 53.150 147.610 53.350 ;
        RECT 147.315 51.750 147.775 53.150 ;
        RECT 146.705 49.550 147.165 50.950 ;
        RECT 146.740 49.350 146.970 49.550 ;
        RECT 147.380 49.350 147.610 51.750 ;
        RECT 148.020 50.950 148.250 53.350 ;
        RECT 147.990 49.550 148.350 50.950 ;
        RECT 148.020 49.350 148.250 49.550 ;
        RECT 148.970 49.200 149.240 53.500 ;
        RECT 135.140 48.900 143.240 49.200 ;
        RECT 145.090 48.900 149.240 49.200 ;
        RECT 16.600 46.680 21.760 46.910 ;
        RECT 16.600 46.660 21.735 46.680 ;
        RECT 16.600 46.610 17.050 46.660 ;
        RECT 24.025 46.595 24.475 46.915 ;
        RECT 10.250 38.495 10.600 46.485 ;
        RECT 11.600 45.585 19.700 45.885 ;
        RECT 11.320 43.160 11.550 45.405 ;
        RECT 11.275 41.760 11.735 43.160 ;
        RECT 11.320 39.405 11.550 41.760 ;
        RECT 11.960 40.960 12.190 45.405 ;
        RECT 12.600 43.160 12.830 45.405 ;
        RECT 12.550 41.760 13.010 43.160 ;
        RECT 11.925 39.560 12.385 40.960 ;
        RECT 11.960 39.405 12.190 39.560 ;
        RECT 12.600 39.405 12.830 41.760 ;
        RECT 13.240 40.960 13.470 45.405 ;
        RECT 13.880 43.160 14.110 45.405 ;
        RECT 13.825 41.760 14.285 43.160 ;
        RECT 13.215 39.560 13.675 40.960 ;
        RECT 13.240 39.405 13.470 39.560 ;
        RECT 13.880 39.405 14.110 41.760 ;
        RECT 14.520 40.960 14.750 45.405 ;
        RECT 15.160 43.160 15.390 45.405 ;
        RECT 15.100 41.760 15.560 43.160 ;
        RECT 14.490 39.560 14.950 40.960 ;
        RECT 14.520 39.405 14.750 39.560 ;
        RECT 15.160 39.405 15.390 41.760 ;
        RECT 15.800 40.960 16.030 45.405 ;
        RECT 16.440 43.160 16.670 45.405 ;
        RECT 16.375 41.760 16.835 43.160 ;
        RECT 15.765 39.560 16.225 40.960 ;
        RECT 15.800 39.405 16.030 39.560 ;
        RECT 16.440 39.405 16.670 41.760 ;
        RECT 17.080 40.960 17.310 45.405 ;
        RECT 17.720 43.160 17.950 45.405 ;
        RECT 17.650 41.760 18.110 43.160 ;
        RECT 17.040 39.560 17.500 40.960 ;
        RECT 17.080 39.405 17.310 39.560 ;
        RECT 17.720 39.405 17.950 41.760 ;
        RECT 18.360 40.960 18.590 45.405 ;
        RECT 19.300 44.410 19.700 45.585 ;
        RECT 25.350 44.410 25.700 44.460 ;
        RECT 19.300 44.110 25.700 44.410 ;
        RECT 18.315 39.560 18.775 40.960 ;
        RECT 18.360 39.405 18.590 39.560 ;
        RECT 19.300 39.210 19.700 44.110 ;
        RECT 25.350 44.060 25.700 44.110 ;
        RECT 21.550 43.510 25.700 43.810 ;
        RECT 21.280 43.160 21.510 43.360 ;
        RECT 21.225 41.760 21.685 43.160 ;
        RECT 21.280 39.360 21.510 41.760 ;
        RECT 21.920 40.960 22.150 43.360 ;
        RECT 22.560 43.160 22.790 43.360 ;
        RECT 22.500 41.760 22.960 43.160 ;
        RECT 21.890 39.560 22.350 40.960 ;
        RECT 21.920 39.360 22.150 39.560 ;
        RECT 22.560 39.360 22.790 41.760 ;
        RECT 23.200 40.960 23.430 43.360 ;
        RECT 23.840 43.160 24.070 43.360 ;
        RECT 23.775 41.760 24.235 43.160 ;
        RECT 23.165 39.560 23.625 40.960 ;
        RECT 23.200 39.360 23.430 39.560 ;
        RECT 23.840 39.360 24.070 41.760 ;
        RECT 24.480 40.960 24.710 43.360 ;
        RECT 25.430 42.760 25.700 43.510 ;
        RECT 25.350 42.360 25.700 42.760 ;
        RECT 24.450 39.560 24.810 40.960 ;
        RECT 24.480 39.360 24.710 39.560 ;
        RECT 25.430 39.210 25.700 42.360 ;
        RECT 11.600 38.910 19.700 39.210 ;
        RECT 8.050 37.430 17.300 38.495 ;
        RECT 17.920 38.010 18.150 38.100 ;
        RECT 18.360 38.010 18.590 38.100 ;
        RECT 19.300 38.010 19.700 38.910 ;
        RECT 20.160 38.910 25.700 39.210 ;
        RECT 17.815 37.660 18.175 38.010 ;
        RECT 18.340 37.660 18.700 38.010 ;
        RECT 19.250 37.660 19.750 38.010 ;
        RECT 17.920 37.100 18.150 37.660 ;
        RECT 18.360 37.100 18.590 37.660 ;
        RECT 19.300 37.610 19.700 37.660 ;
        RECT 16.600 36.910 17.050 36.960 ;
        RECT 20.160 36.910 20.560 38.910 ;
        RECT 25.850 38.760 26.200 47.430 ;
        RECT 133.655 47.420 140.840 48.485 ;
        RECT 141.460 48.000 141.690 48.090 ;
        RECT 141.900 48.000 142.130 48.090 ;
        RECT 142.840 48.000 143.240 48.900 ;
        RECT 144.820 48.000 145.050 48.060 ;
        RECT 145.260 48.000 145.490 48.060 ;
        RECT 141.355 47.650 141.715 48.000 ;
        RECT 141.880 47.650 142.240 48.000 ;
        RECT 142.790 47.650 143.290 48.000 ;
        RECT 144.705 47.650 145.065 48.000 ;
        RECT 145.230 47.650 145.590 48.000 ;
        RECT 141.460 47.090 141.690 47.650 ;
        RECT 141.900 47.090 142.130 47.650 ;
        RECT 142.840 47.600 143.240 47.650 ;
        RECT 144.820 47.060 145.050 47.650 ;
        RECT 145.260 47.060 145.490 47.650 ;
        RECT 146.390 46.955 146.690 48.900 ;
        RECT 149.390 48.485 149.740 56.475 ;
        RECT 146.840 47.420 151.990 48.485 ;
        RECT 139.690 46.900 140.090 46.950 ;
        RECT 146.335 46.900 146.745 46.955 ;
        RECT 139.690 46.650 146.745 46.900 ;
        RECT 139.690 46.600 140.090 46.650 ;
        RECT 146.335 46.595 146.745 46.650 ;
        RECT 22.670 38.560 26.200 38.760 ;
        RECT 21.280 38.010 21.510 38.070 ;
        RECT 21.720 38.010 21.950 38.070 ;
        RECT 21.165 37.660 21.525 38.010 ;
        RECT 21.690 37.660 22.050 38.010 ;
        RECT 22.670 37.660 23.200 38.560 ;
        RECT 25.100 38.495 26.200 38.560 ;
        RECT 23.920 38.010 24.150 38.060 ;
        RECT 23.775 37.660 24.150 38.010 ;
        RECT 21.280 37.070 21.510 37.660 ;
        RECT 21.720 37.070 21.950 37.660 ;
        RECT 23.920 37.060 24.150 37.660 ;
        RECT 24.360 38.010 24.590 38.060 ;
        RECT 24.360 37.660 24.740 38.010 ;
        RECT 24.360 37.060 24.590 37.660 ;
        RECT 25.100 37.430 26.335 38.495 ;
        RECT 133.790 38.485 134.140 46.475 ;
        RECT 134.290 45.875 134.640 45.925 ;
        RECT 134.290 45.575 143.240 45.875 ;
        RECT 134.860 43.150 135.090 45.395 ;
        RECT 134.815 41.750 135.275 43.150 ;
        RECT 134.860 39.395 135.090 41.750 ;
        RECT 135.500 40.950 135.730 45.395 ;
        RECT 136.140 43.150 136.370 45.395 ;
        RECT 136.090 41.750 136.550 43.150 ;
        RECT 135.465 39.550 135.925 40.950 ;
        RECT 135.500 39.395 135.730 39.550 ;
        RECT 136.140 39.395 136.370 41.750 ;
        RECT 136.780 40.950 137.010 45.395 ;
        RECT 137.420 43.150 137.650 45.395 ;
        RECT 137.365 41.750 137.825 43.150 ;
        RECT 136.755 39.550 137.215 40.950 ;
        RECT 136.780 39.395 137.010 39.550 ;
        RECT 137.420 39.395 137.650 41.750 ;
        RECT 138.060 40.950 138.290 45.395 ;
        RECT 138.700 43.150 138.930 45.395 ;
        RECT 138.640 41.750 139.100 43.150 ;
        RECT 138.030 39.550 138.490 40.950 ;
        RECT 138.060 39.395 138.290 39.550 ;
        RECT 138.700 39.395 138.930 41.750 ;
        RECT 139.340 40.950 139.570 45.395 ;
        RECT 139.980 43.150 140.210 45.395 ;
        RECT 139.915 41.750 140.375 43.150 ;
        RECT 139.305 39.550 139.765 40.950 ;
        RECT 139.340 39.395 139.570 39.550 ;
        RECT 139.980 39.395 140.210 41.750 ;
        RECT 140.620 40.950 140.850 45.395 ;
        RECT 141.260 43.150 141.490 45.395 ;
        RECT 141.190 41.750 141.650 43.150 ;
        RECT 140.580 39.550 141.040 40.950 ;
        RECT 140.620 39.395 140.850 39.550 ;
        RECT 141.260 39.395 141.490 41.750 ;
        RECT 141.900 40.950 142.130 45.395 ;
        RECT 141.855 39.550 142.315 40.950 ;
        RECT 141.900 39.395 142.130 39.550 ;
        RECT 142.840 39.200 143.240 45.575 ;
        RECT 145.090 43.500 149.240 43.800 ;
        RECT 144.820 43.150 145.050 43.350 ;
        RECT 144.765 41.750 145.225 43.150 ;
        RECT 144.820 39.350 145.050 41.750 ;
        RECT 145.460 40.950 145.690 43.350 ;
        RECT 146.100 43.150 146.330 43.350 ;
        RECT 146.040 41.750 146.500 43.150 ;
        RECT 145.430 39.550 145.890 40.950 ;
        RECT 145.460 39.350 145.690 39.550 ;
        RECT 146.100 39.350 146.330 41.750 ;
        RECT 146.740 40.950 146.970 43.350 ;
        RECT 147.380 43.150 147.610 43.350 ;
        RECT 147.315 41.750 147.775 43.150 ;
        RECT 146.705 39.550 147.165 40.950 ;
        RECT 146.740 39.350 146.970 39.550 ;
        RECT 147.380 39.350 147.610 41.750 ;
        RECT 148.020 40.950 148.250 43.350 ;
        RECT 147.990 39.550 148.350 40.950 ;
        RECT 148.020 39.350 148.250 39.550 ;
        RECT 148.970 39.200 149.240 43.500 ;
        RECT 135.140 38.900 143.240 39.200 ;
        RECT 145.090 38.900 149.240 39.200 ;
        RECT 16.600 36.680 21.760 36.910 ;
        RECT 16.600 36.660 21.735 36.680 ;
        RECT 16.600 36.610 17.050 36.660 ;
        RECT 24.025 36.595 24.475 36.915 ;
        RECT 10.250 28.495 10.600 36.485 ;
        RECT 11.600 35.585 19.700 35.885 ;
        RECT 11.320 33.160 11.550 35.405 ;
        RECT 11.275 31.760 11.735 33.160 ;
        RECT 11.320 29.405 11.550 31.760 ;
        RECT 11.960 30.960 12.190 35.405 ;
        RECT 12.600 33.160 12.830 35.405 ;
        RECT 12.550 31.760 13.010 33.160 ;
        RECT 11.925 29.560 12.385 30.960 ;
        RECT 11.960 29.405 12.190 29.560 ;
        RECT 12.600 29.405 12.830 31.760 ;
        RECT 13.240 30.960 13.470 35.405 ;
        RECT 13.880 33.160 14.110 35.405 ;
        RECT 13.825 31.760 14.285 33.160 ;
        RECT 13.215 29.560 13.675 30.960 ;
        RECT 13.240 29.405 13.470 29.560 ;
        RECT 13.880 29.405 14.110 31.760 ;
        RECT 14.520 30.960 14.750 35.405 ;
        RECT 15.160 33.160 15.390 35.405 ;
        RECT 15.100 31.760 15.560 33.160 ;
        RECT 14.490 29.560 14.950 30.960 ;
        RECT 14.520 29.405 14.750 29.560 ;
        RECT 15.160 29.405 15.390 31.760 ;
        RECT 15.800 30.960 16.030 35.405 ;
        RECT 16.440 33.160 16.670 35.405 ;
        RECT 16.375 31.760 16.835 33.160 ;
        RECT 15.765 29.560 16.225 30.960 ;
        RECT 15.800 29.405 16.030 29.560 ;
        RECT 16.440 29.405 16.670 31.760 ;
        RECT 17.080 30.960 17.310 35.405 ;
        RECT 17.720 33.160 17.950 35.405 ;
        RECT 17.650 31.760 18.110 33.160 ;
        RECT 17.040 29.560 17.500 30.960 ;
        RECT 17.080 29.405 17.310 29.560 ;
        RECT 17.720 29.405 17.950 31.760 ;
        RECT 18.360 30.960 18.590 35.405 ;
        RECT 19.300 34.410 19.700 35.585 ;
        RECT 25.350 34.410 25.700 34.460 ;
        RECT 19.300 34.110 25.700 34.410 ;
        RECT 18.315 29.560 18.775 30.960 ;
        RECT 18.360 29.405 18.590 29.560 ;
        RECT 19.300 29.210 19.700 34.110 ;
        RECT 25.350 34.060 25.700 34.110 ;
        RECT 21.550 33.510 25.700 33.810 ;
        RECT 21.280 33.160 21.510 33.360 ;
        RECT 21.225 31.760 21.685 33.160 ;
        RECT 21.280 29.360 21.510 31.760 ;
        RECT 21.920 30.960 22.150 33.360 ;
        RECT 22.560 33.160 22.790 33.360 ;
        RECT 22.500 31.760 22.960 33.160 ;
        RECT 21.890 29.560 22.350 30.960 ;
        RECT 21.920 29.360 22.150 29.560 ;
        RECT 22.560 29.360 22.790 31.760 ;
        RECT 23.200 30.960 23.430 33.360 ;
        RECT 23.840 33.160 24.070 33.360 ;
        RECT 23.775 31.760 24.235 33.160 ;
        RECT 23.165 29.560 23.625 30.960 ;
        RECT 23.200 29.360 23.430 29.560 ;
        RECT 23.840 29.360 24.070 31.760 ;
        RECT 24.480 30.960 24.710 33.360 ;
        RECT 25.430 32.760 25.700 33.510 ;
        RECT 25.350 32.360 25.700 32.760 ;
        RECT 24.450 29.560 24.810 30.960 ;
        RECT 24.480 29.360 24.710 29.560 ;
        RECT 25.430 29.210 25.700 32.360 ;
        RECT 11.600 28.910 19.700 29.210 ;
        RECT 8.050 27.430 17.300 28.495 ;
        RECT 17.920 28.010 18.150 28.100 ;
        RECT 18.360 28.010 18.590 28.100 ;
        RECT 19.300 28.010 19.700 28.910 ;
        RECT 20.160 28.910 25.700 29.210 ;
        RECT 17.815 27.660 18.175 28.010 ;
        RECT 18.340 27.660 18.700 28.010 ;
        RECT 19.250 27.660 19.750 28.010 ;
        RECT 17.920 27.100 18.150 27.660 ;
        RECT 18.360 27.100 18.590 27.660 ;
        RECT 19.300 27.610 19.700 27.660 ;
        RECT 16.600 26.910 17.050 26.960 ;
        RECT 20.160 26.910 20.560 28.910 ;
        RECT 25.850 28.760 26.200 37.430 ;
        RECT 133.655 37.420 140.840 38.485 ;
        RECT 141.460 38.000 141.690 38.090 ;
        RECT 141.900 38.000 142.130 38.090 ;
        RECT 142.840 38.000 143.240 38.900 ;
        RECT 144.820 38.000 145.050 38.060 ;
        RECT 145.260 38.000 145.490 38.060 ;
        RECT 141.355 37.650 141.715 38.000 ;
        RECT 141.880 37.650 142.240 38.000 ;
        RECT 142.790 37.650 143.290 38.000 ;
        RECT 144.705 37.650 145.065 38.000 ;
        RECT 145.230 37.650 145.590 38.000 ;
        RECT 141.460 37.090 141.690 37.650 ;
        RECT 141.900 37.090 142.130 37.650 ;
        RECT 142.840 37.600 143.240 37.650 ;
        RECT 144.820 37.060 145.050 37.650 ;
        RECT 145.260 37.060 145.490 37.650 ;
        RECT 146.390 36.955 146.690 38.900 ;
        RECT 149.390 38.485 149.740 46.475 ;
        RECT 146.840 37.420 151.990 38.485 ;
        RECT 139.690 36.900 140.090 36.950 ;
        RECT 146.335 36.900 146.745 36.955 ;
        RECT 139.690 36.650 146.745 36.900 ;
        RECT 139.690 36.600 140.090 36.650 ;
        RECT 146.335 36.595 146.745 36.650 ;
        RECT 22.670 28.560 26.200 28.760 ;
        RECT 21.280 28.010 21.510 28.070 ;
        RECT 21.720 28.010 21.950 28.070 ;
        RECT 21.165 27.660 21.525 28.010 ;
        RECT 21.690 27.660 22.050 28.010 ;
        RECT 22.670 27.660 23.200 28.560 ;
        RECT 25.100 28.495 26.200 28.560 ;
        RECT 23.920 28.010 24.150 28.060 ;
        RECT 23.775 27.660 24.150 28.010 ;
        RECT 21.280 27.070 21.510 27.660 ;
        RECT 21.720 27.070 21.950 27.660 ;
        RECT 23.920 27.060 24.150 27.660 ;
        RECT 24.360 28.010 24.590 28.060 ;
        RECT 24.360 27.660 24.740 28.010 ;
        RECT 24.360 27.060 24.590 27.660 ;
        RECT 25.100 27.430 26.335 28.495 ;
        RECT 133.790 28.485 134.140 36.475 ;
        RECT 134.290 35.875 134.640 35.925 ;
        RECT 134.290 35.575 143.240 35.875 ;
        RECT 134.860 33.150 135.090 35.395 ;
        RECT 134.815 31.750 135.275 33.150 ;
        RECT 134.860 29.395 135.090 31.750 ;
        RECT 135.500 30.950 135.730 35.395 ;
        RECT 136.140 33.150 136.370 35.395 ;
        RECT 136.090 31.750 136.550 33.150 ;
        RECT 135.465 29.550 135.925 30.950 ;
        RECT 135.500 29.395 135.730 29.550 ;
        RECT 136.140 29.395 136.370 31.750 ;
        RECT 136.780 30.950 137.010 35.395 ;
        RECT 137.420 33.150 137.650 35.395 ;
        RECT 137.365 31.750 137.825 33.150 ;
        RECT 136.755 29.550 137.215 30.950 ;
        RECT 136.780 29.395 137.010 29.550 ;
        RECT 137.420 29.395 137.650 31.750 ;
        RECT 138.060 30.950 138.290 35.395 ;
        RECT 138.700 33.150 138.930 35.395 ;
        RECT 138.640 31.750 139.100 33.150 ;
        RECT 138.030 29.550 138.490 30.950 ;
        RECT 138.060 29.395 138.290 29.550 ;
        RECT 138.700 29.395 138.930 31.750 ;
        RECT 139.340 30.950 139.570 35.395 ;
        RECT 139.980 33.150 140.210 35.395 ;
        RECT 139.915 31.750 140.375 33.150 ;
        RECT 139.305 29.550 139.765 30.950 ;
        RECT 139.340 29.395 139.570 29.550 ;
        RECT 139.980 29.395 140.210 31.750 ;
        RECT 140.620 30.950 140.850 35.395 ;
        RECT 141.260 33.150 141.490 35.395 ;
        RECT 141.190 31.750 141.650 33.150 ;
        RECT 140.580 29.550 141.040 30.950 ;
        RECT 140.620 29.395 140.850 29.550 ;
        RECT 141.260 29.395 141.490 31.750 ;
        RECT 141.900 30.950 142.130 35.395 ;
        RECT 141.855 29.550 142.315 30.950 ;
        RECT 141.900 29.395 142.130 29.550 ;
        RECT 142.840 29.200 143.240 35.575 ;
        RECT 145.090 33.500 149.240 33.800 ;
        RECT 144.820 33.150 145.050 33.350 ;
        RECT 144.765 31.750 145.225 33.150 ;
        RECT 144.820 29.350 145.050 31.750 ;
        RECT 145.460 30.950 145.690 33.350 ;
        RECT 146.100 33.150 146.330 33.350 ;
        RECT 146.040 31.750 146.500 33.150 ;
        RECT 145.430 29.550 145.890 30.950 ;
        RECT 145.460 29.350 145.690 29.550 ;
        RECT 146.100 29.350 146.330 31.750 ;
        RECT 146.740 30.950 146.970 33.350 ;
        RECT 147.380 33.150 147.610 33.350 ;
        RECT 147.315 31.750 147.775 33.150 ;
        RECT 146.705 29.550 147.165 30.950 ;
        RECT 146.740 29.350 146.970 29.550 ;
        RECT 147.380 29.350 147.610 31.750 ;
        RECT 148.020 30.950 148.250 33.350 ;
        RECT 147.990 29.550 148.350 30.950 ;
        RECT 148.020 29.350 148.250 29.550 ;
        RECT 148.970 29.200 149.240 33.500 ;
        RECT 135.140 28.900 143.240 29.200 ;
        RECT 145.090 28.900 149.240 29.200 ;
        RECT 16.600 26.680 21.760 26.910 ;
        RECT 16.600 26.660 21.735 26.680 ;
        RECT 16.600 26.610 17.050 26.660 ;
        RECT 24.025 26.595 24.475 26.915 ;
        RECT 10.250 18.495 10.600 26.485 ;
        RECT 11.600 25.585 19.700 25.885 ;
        RECT 11.320 23.160 11.550 25.405 ;
        RECT 11.275 21.760 11.735 23.160 ;
        RECT 11.320 19.405 11.550 21.760 ;
        RECT 11.960 20.960 12.190 25.405 ;
        RECT 12.600 23.160 12.830 25.405 ;
        RECT 12.550 21.760 13.010 23.160 ;
        RECT 11.925 19.560 12.385 20.960 ;
        RECT 11.960 19.405 12.190 19.560 ;
        RECT 12.600 19.405 12.830 21.760 ;
        RECT 13.240 20.960 13.470 25.405 ;
        RECT 13.880 23.160 14.110 25.405 ;
        RECT 13.825 21.760 14.285 23.160 ;
        RECT 13.215 19.560 13.675 20.960 ;
        RECT 13.240 19.405 13.470 19.560 ;
        RECT 13.880 19.405 14.110 21.760 ;
        RECT 14.520 20.960 14.750 25.405 ;
        RECT 15.160 23.160 15.390 25.405 ;
        RECT 15.100 21.760 15.560 23.160 ;
        RECT 14.490 19.560 14.950 20.960 ;
        RECT 14.520 19.405 14.750 19.560 ;
        RECT 15.160 19.405 15.390 21.760 ;
        RECT 15.800 20.960 16.030 25.405 ;
        RECT 16.440 23.160 16.670 25.405 ;
        RECT 16.375 21.760 16.835 23.160 ;
        RECT 15.765 19.560 16.225 20.960 ;
        RECT 15.800 19.405 16.030 19.560 ;
        RECT 16.440 19.405 16.670 21.760 ;
        RECT 17.080 20.960 17.310 25.405 ;
        RECT 17.720 23.160 17.950 25.405 ;
        RECT 17.650 21.760 18.110 23.160 ;
        RECT 17.040 19.560 17.500 20.960 ;
        RECT 17.080 19.405 17.310 19.560 ;
        RECT 17.720 19.405 17.950 21.760 ;
        RECT 18.360 20.960 18.590 25.405 ;
        RECT 19.300 24.410 19.700 25.585 ;
        RECT 25.350 24.410 25.700 24.460 ;
        RECT 19.300 24.110 25.700 24.410 ;
        RECT 18.315 19.560 18.775 20.960 ;
        RECT 18.360 19.405 18.590 19.560 ;
        RECT 19.300 19.210 19.700 24.110 ;
        RECT 25.350 24.060 25.700 24.110 ;
        RECT 21.550 23.510 25.700 23.810 ;
        RECT 21.280 23.160 21.510 23.360 ;
        RECT 21.225 21.760 21.685 23.160 ;
        RECT 21.280 19.360 21.510 21.760 ;
        RECT 21.920 20.960 22.150 23.360 ;
        RECT 22.560 23.160 22.790 23.360 ;
        RECT 22.500 21.760 22.960 23.160 ;
        RECT 21.890 19.560 22.350 20.960 ;
        RECT 21.920 19.360 22.150 19.560 ;
        RECT 22.560 19.360 22.790 21.760 ;
        RECT 23.200 20.960 23.430 23.360 ;
        RECT 23.840 23.160 24.070 23.360 ;
        RECT 23.775 21.760 24.235 23.160 ;
        RECT 23.165 19.560 23.625 20.960 ;
        RECT 23.200 19.360 23.430 19.560 ;
        RECT 23.840 19.360 24.070 21.760 ;
        RECT 24.480 20.960 24.710 23.360 ;
        RECT 25.430 22.760 25.700 23.510 ;
        RECT 25.350 22.360 25.700 22.760 ;
        RECT 24.450 19.560 24.810 20.960 ;
        RECT 24.480 19.360 24.710 19.560 ;
        RECT 25.430 19.210 25.700 22.360 ;
        RECT 11.600 18.910 19.700 19.210 ;
        RECT 8.050 17.430 17.300 18.495 ;
        RECT 17.920 18.010 18.150 18.100 ;
        RECT 18.360 18.010 18.590 18.100 ;
        RECT 19.300 18.010 19.700 18.910 ;
        RECT 20.160 18.910 25.700 19.210 ;
        RECT 17.815 17.660 18.175 18.010 ;
        RECT 18.340 17.660 18.700 18.010 ;
        RECT 19.250 17.660 19.750 18.010 ;
        RECT 17.920 17.100 18.150 17.660 ;
        RECT 18.360 17.100 18.590 17.660 ;
        RECT 19.300 17.610 19.700 17.660 ;
        RECT 16.600 16.910 17.050 16.960 ;
        RECT 20.160 16.910 20.560 18.910 ;
        RECT 25.850 18.760 26.200 27.430 ;
        RECT 133.655 27.420 140.840 28.485 ;
        RECT 141.460 28.000 141.690 28.090 ;
        RECT 141.900 28.000 142.130 28.090 ;
        RECT 142.840 28.000 143.240 28.900 ;
        RECT 144.820 28.000 145.050 28.060 ;
        RECT 145.260 28.000 145.490 28.060 ;
        RECT 141.355 27.650 141.715 28.000 ;
        RECT 141.880 27.650 142.240 28.000 ;
        RECT 142.790 27.650 143.290 28.000 ;
        RECT 144.705 27.650 145.065 28.000 ;
        RECT 145.230 27.650 145.590 28.000 ;
        RECT 141.460 27.090 141.690 27.650 ;
        RECT 141.900 27.090 142.130 27.650 ;
        RECT 142.840 27.600 143.240 27.650 ;
        RECT 144.820 27.060 145.050 27.650 ;
        RECT 145.260 27.060 145.490 27.650 ;
        RECT 146.390 26.955 146.690 28.900 ;
        RECT 149.390 28.485 149.740 36.475 ;
        RECT 146.840 27.420 151.990 28.485 ;
        RECT 139.690 26.900 140.090 26.950 ;
        RECT 146.335 26.900 146.745 26.955 ;
        RECT 139.690 26.650 146.745 26.900 ;
        RECT 139.690 26.600 140.090 26.650 ;
        RECT 146.335 26.595 146.745 26.650 ;
        RECT 22.670 18.560 26.200 18.760 ;
        RECT 21.280 18.010 21.510 18.070 ;
        RECT 21.720 18.010 21.950 18.070 ;
        RECT 21.165 17.660 21.525 18.010 ;
        RECT 21.690 17.660 22.050 18.010 ;
        RECT 22.670 17.660 23.200 18.560 ;
        RECT 25.100 18.495 26.200 18.560 ;
        RECT 23.920 18.010 24.150 18.060 ;
        RECT 23.775 17.660 24.150 18.010 ;
        RECT 21.280 17.070 21.510 17.660 ;
        RECT 21.720 17.070 21.950 17.660 ;
        RECT 23.920 17.060 24.150 17.660 ;
        RECT 24.360 18.010 24.590 18.060 ;
        RECT 24.360 17.660 24.740 18.010 ;
        RECT 24.360 17.060 24.590 17.660 ;
        RECT 25.100 17.430 26.335 18.495 ;
        RECT 133.790 18.485 134.140 26.475 ;
        RECT 134.290 25.875 134.640 25.925 ;
        RECT 134.290 25.575 143.240 25.875 ;
        RECT 134.860 23.150 135.090 25.395 ;
        RECT 134.815 21.750 135.275 23.150 ;
        RECT 134.860 19.395 135.090 21.750 ;
        RECT 135.500 20.950 135.730 25.395 ;
        RECT 136.140 23.150 136.370 25.395 ;
        RECT 136.090 21.750 136.550 23.150 ;
        RECT 135.465 19.550 135.925 20.950 ;
        RECT 135.500 19.395 135.730 19.550 ;
        RECT 136.140 19.395 136.370 21.750 ;
        RECT 136.780 20.950 137.010 25.395 ;
        RECT 137.420 23.150 137.650 25.395 ;
        RECT 137.365 21.750 137.825 23.150 ;
        RECT 136.755 19.550 137.215 20.950 ;
        RECT 136.780 19.395 137.010 19.550 ;
        RECT 137.420 19.395 137.650 21.750 ;
        RECT 138.060 20.950 138.290 25.395 ;
        RECT 138.700 23.150 138.930 25.395 ;
        RECT 138.640 21.750 139.100 23.150 ;
        RECT 138.030 19.550 138.490 20.950 ;
        RECT 138.060 19.395 138.290 19.550 ;
        RECT 138.700 19.395 138.930 21.750 ;
        RECT 139.340 20.950 139.570 25.395 ;
        RECT 139.980 23.150 140.210 25.395 ;
        RECT 139.915 21.750 140.375 23.150 ;
        RECT 139.305 19.550 139.765 20.950 ;
        RECT 139.340 19.395 139.570 19.550 ;
        RECT 139.980 19.395 140.210 21.750 ;
        RECT 140.620 20.950 140.850 25.395 ;
        RECT 141.260 23.150 141.490 25.395 ;
        RECT 141.190 21.750 141.650 23.150 ;
        RECT 140.580 19.550 141.040 20.950 ;
        RECT 140.620 19.395 140.850 19.550 ;
        RECT 141.260 19.395 141.490 21.750 ;
        RECT 141.900 20.950 142.130 25.395 ;
        RECT 141.855 19.550 142.315 20.950 ;
        RECT 141.900 19.395 142.130 19.550 ;
        RECT 142.840 19.200 143.240 25.575 ;
        RECT 145.090 23.500 149.240 23.800 ;
        RECT 144.820 23.150 145.050 23.350 ;
        RECT 144.765 21.750 145.225 23.150 ;
        RECT 144.820 19.350 145.050 21.750 ;
        RECT 145.460 20.950 145.690 23.350 ;
        RECT 146.100 23.150 146.330 23.350 ;
        RECT 146.040 21.750 146.500 23.150 ;
        RECT 145.430 19.550 145.890 20.950 ;
        RECT 145.460 19.350 145.690 19.550 ;
        RECT 146.100 19.350 146.330 21.750 ;
        RECT 146.740 20.950 146.970 23.350 ;
        RECT 147.380 23.150 147.610 23.350 ;
        RECT 147.315 21.750 147.775 23.150 ;
        RECT 146.705 19.550 147.165 20.950 ;
        RECT 146.740 19.350 146.970 19.550 ;
        RECT 147.380 19.350 147.610 21.750 ;
        RECT 148.020 20.950 148.250 23.350 ;
        RECT 147.990 19.550 148.350 20.950 ;
        RECT 148.020 19.350 148.250 19.550 ;
        RECT 148.970 19.200 149.240 23.500 ;
        RECT 135.140 18.900 143.240 19.200 ;
        RECT 145.090 18.900 149.240 19.200 ;
        RECT 16.600 16.680 21.760 16.910 ;
        RECT 16.600 16.660 21.735 16.680 ;
        RECT 16.600 16.610 17.050 16.660 ;
        RECT 24.025 16.595 24.475 16.915 ;
        RECT 10.250 8.495 10.600 16.485 ;
        RECT 11.600 15.585 19.700 15.885 ;
        RECT 11.320 13.160 11.550 15.405 ;
        RECT 11.275 11.760 11.735 13.160 ;
        RECT 11.320 9.405 11.550 11.760 ;
        RECT 11.960 10.960 12.190 15.405 ;
        RECT 12.600 13.160 12.830 15.405 ;
        RECT 12.550 11.760 13.010 13.160 ;
        RECT 11.925 9.560 12.385 10.960 ;
        RECT 11.960 9.405 12.190 9.560 ;
        RECT 12.600 9.405 12.830 11.760 ;
        RECT 13.240 10.960 13.470 15.405 ;
        RECT 13.880 13.160 14.110 15.405 ;
        RECT 13.825 11.760 14.285 13.160 ;
        RECT 13.215 9.560 13.675 10.960 ;
        RECT 13.240 9.405 13.470 9.560 ;
        RECT 13.880 9.405 14.110 11.760 ;
        RECT 14.520 10.960 14.750 15.405 ;
        RECT 15.160 13.160 15.390 15.405 ;
        RECT 15.100 11.760 15.560 13.160 ;
        RECT 14.490 9.560 14.950 10.960 ;
        RECT 14.520 9.405 14.750 9.560 ;
        RECT 15.160 9.405 15.390 11.760 ;
        RECT 15.800 10.960 16.030 15.405 ;
        RECT 16.440 13.160 16.670 15.405 ;
        RECT 16.375 11.760 16.835 13.160 ;
        RECT 15.765 9.560 16.225 10.960 ;
        RECT 15.800 9.405 16.030 9.560 ;
        RECT 16.440 9.405 16.670 11.760 ;
        RECT 17.080 10.960 17.310 15.405 ;
        RECT 17.720 13.160 17.950 15.405 ;
        RECT 17.650 11.760 18.110 13.160 ;
        RECT 17.040 9.560 17.500 10.960 ;
        RECT 17.080 9.405 17.310 9.560 ;
        RECT 17.720 9.405 17.950 11.760 ;
        RECT 18.360 10.960 18.590 15.405 ;
        RECT 19.300 14.410 19.700 15.585 ;
        RECT 25.350 14.410 25.700 14.460 ;
        RECT 19.300 14.110 25.700 14.410 ;
        RECT 18.315 9.560 18.775 10.960 ;
        RECT 18.360 9.405 18.590 9.560 ;
        RECT 19.300 9.210 19.700 14.110 ;
        RECT 25.350 14.060 25.700 14.110 ;
        RECT 21.550 13.510 25.700 13.810 ;
        RECT 21.280 13.160 21.510 13.360 ;
        RECT 21.225 11.760 21.685 13.160 ;
        RECT 21.280 9.360 21.510 11.760 ;
        RECT 21.920 10.960 22.150 13.360 ;
        RECT 22.560 13.160 22.790 13.360 ;
        RECT 22.500 11.760 22.960 13.160 ;
        RECT 21.890 9.560 22.350 10.960 ;
        RECT 21.920 9.360 22.150 9.560 ;
        RECT 22.560 9.360 22.790 11.760 ;
        RECT 23.200 10.960 23.430 13.360 ;
        RECT 23.840 13.160 24.070 13.360 ;
        RECT 23.775 11.760 24.235 13.160 ;
        RECT 23.165 9.560 23.625 10.960 ;
        RECT 23.200 9.360 23.430 9.560 ;
        RECT 23.840 9.360 24.070 11.760 ;
        RECT 24.480 10.960 24.710 13.360 ;
        RECT 25.430 12.760 25.700 13.510 ;
        RECT 25.350 12.360 25.700 12.760 ;
        RECT 24.450 9.560 24.810 10.960 ;
        RECT 24.480 9.360 24.710 9.560 ;
        RECT 25.430 9.210 25.700 12.360 ;
        RECT 11.600 8.910 19.700 9.210 ;
        RECT 8.050 7.430 17.300 8.495 ;
        RECT 17.920 8.010 18.150 8.100 ;
        RECT 18.360 8.010 18.590 8.100 ;
        RECT 19.300 8.010 19.700 8.910 ;
        RECT 20.160 8.910 25.700 9.210 ;
        RECT 17.815 7.660 18.175 8.010 ;
        RECT 18.340 7.660 18.700 8.010 ;
        RECT 19.250 7.660 19.750 8.010 ;
        RECT 17.920 7.100 18.150 7.660 ;
        RECT 18.360 7.100 18.590 7.660 ;
        RECT 19.300 7.610 19.700 7.660 ;
        RECT 16.600 6.910 17.050 6.960 ;
        RECT 20.160 6.910 20.560 8.910 ;
        RECT 25.850 8.760 26.200 17.430 ;
        RECT 133.655 17.420 140.840 18.485 ;
        RECT 141.460 18.000 141.690 18.090 ;
        RECT 141.900 18.000 142.130 18.090 ;
        RECT 142.840 18.000 143.240 18.900 ;
        RECT 144.820 18.000 145.050 18.060 ;
        RECT 145.260 18.000 145.490 18.060 ;
        RECT 141.355 17.650 141.715 18.000 ;
        RECT 141.880 17.650 142.240 18.000 ;
        RECT 142.790 17.650 143.290 18.000 ;
        RECT 144.705 17.650 145.065 18.000 ;
        RECT 145.230 17.650 145.590 18.000 ;
        RECT 141.460 17.090 141.690 17.650 ;
        RECT 141.900 17.090 142.130 17.650 ;
        RECT 142.840 17.600 143.240 17.650 ;
        RECT 144.820 17.060 145.050 17.650 ;
        RECT 145.260 17.060 145.490 17.650 ;
        RECT 146.390 16.955 146.690 18.900 ;
        RECT 149.390 18.485 149.740 26.475 ;
        RECT 146.840 17.420 151.990 18.485 ;
        RECT 139.690 16.900 140.090 16.950 ;
        RECT 146.335 16.900 146.745 16.955 ;
        RECT 139.690 16.650 146.745 16.900 ;
        RECT 139.690 16.600 140.090 16.650 ;
        RECT 146.335 16.595 146.745 16.650 ;
        RECT 22.670 8.560 26.200 8.760 ;
        RECT 21.280 8.010 21.510 8.070 ;
        RECT 21.720 8.010 21.950 8.070 ;
        RECT 21.165 7.660 21.525 8.010 ;
        RECT 21.690 7.660 22.050 8.010 ;
        RECT 22.670 7.660 23.200 8.560 ;
        RECT 25.100 8.495 26.200 8.560 ;
        RECT 23.920 8.010 24.150 8.060 ;
        RECT 23.775 7.660 24.150 8.010 ;
        RECT 21.280 7.070 21.510 7.660 ;
        RECT 21.720 7.070 21.950 7.660 ;
        RECT 23.920 7.060 24.150 7.660 ;
        RECT 24.360 8.010 24.590 8.060 ;
        RECT 24.360 7.660 24.740 8.010 ;
        RECT 24.360 7.060 24.590 7.660 ;
        RECT 25.100 7.430 26.335 8.495 ;
        RECT 133.790 8.485 134.140 16.475 ;
        RECT 134.290 15.875 134.640 15.925 ;
        RECT 134.290 15.575 143.240 15.875 ;
        RECT 134.860 13.150 135.090 15.395 ;
        RECT 134.815 11.750 135.275 13.150 ;
        RECT 134.860 9.395 135.090 11.750 ;
        RECT 135.500 10.950 135.730 15.395 ;
        RECT 136.140 13.150 136.370 15.395 ;
        RECT 136.090 11.750 136.550 13.150 ;
        RECT 135.465 9.550 135.925 10.950 ;
        RECT 135.500 9.395 135.730 9.550 ;
        RECT 136.140 9.395 136.370 11.750 ;
        RECT 136.780 10.950 137.010 15.395 ;
        RECT 137.420 13.150 137.650 15.395 ;
        RECT 137.365 11.750 137.825 13.150 ;
        RECT 136.755 9.550 137.215 10.950 ;
        RECT 136.780 9.395 137.010 9.550 ;
        RECT 137.420 9.395 137.650 11.750 ;
        RECT 138.060 10.950 138.290 15.395 ;
        RECT 138.700 13.150 138.930 15.395 ;
        RECT 138.640 11.750 139.100 13.150 ;
        RECT 138.030 9.550 138.490 10.950 ;
        RECT 138.060 9.395 138.290 9.550 ;
        RECT 138.700 9.395 138.930 11.750 ;
        RECT 139.340 10.950 139.570 15.395 ;
        RECT 139.980 13.150 140.210 15.395 ;
        RECT 139.915 11.750 140.375 13.150 ;
        RECT 139.305 9.550 139.765 10.950 ;
        RECT 139.340 9.395 139.570 9.550 ;
        RECT 139.980 9.395 140.210 11.750 ;
        RECT 140.620 10.950 140.850 15.395 ;
        RECT 141.260 13.150 141.490 15.395 ;
        RECT 141.190 11.750 141.650 13.150 ;
        RECT 140.580 9.550 141.040 10.950 ;
        RECT 140.620 9.395 140.850 9.550 ;
        RECT 141.260 9.395 141.490 11.750 ;
        RECT 141.900 10.950 142.130 15.395 ;
        RECT 141.855 9.550 142.315 10.950 ;
        RECT 141.900 9.395 142.130 9.550 ;
        RECT 142.840 9.200 143.240 15.575 ;
        RECT 145.090 13.500 149.240 13.800 ;
        RECT 144.820 13.150 145.050 13.350 ;
        RECT 144.765 11.750 145.225 13.150 ;
        RECT 144.820 9.350 145.050 11.750 ;
        RECT 145.460 10.950 145.690 13.350 ;
        RECT 146.100 13.150 146.330 13.350 ;
        RECT 146.040 11.750 146.500 13.150 ;
        RECT 145.430 9.550 145.890 10.950 ;
        RECT 145.460 9.350 145.690 9.550 ;
        RECT 146.100 9.350 146.330 11.750 ;
        RECT 146.740 10.950 146.970 13.350 ;
        RECT 147.380 13.150 147.610 13.350 ;
        RECT 147.315 11.750 147.775 13.150 ;
        RECT 146.705 9.550 147.165 10.950 ;
        RECT 146.740 9.350 146.970 9.550 ;
        RECT 147.380 9.350 147.610 11.750 ;
        RECT 148.020 10.950 148.250 13.350 ;
        RECT 147.990 9.550 148.350 10.950 ;
        RECT 148.020 9.350 148.250 9.550 ;
        RECT 148.970 9.200 149.240 13.500 ;
        RECT 135.140 8.900 143.240 9.200 ;
        RECT 145.090 8.900 149.240 9.200 ;
        RECT 16.600 6.680 21.760 6.910 ;
        RECT 16.600 6.660 21.735 6.680 ;
        RECT 16.600 6.610 17.050 6.660 ;
        RECT 24.025 6.595 24.475 6.915 ;
        RECT 25.850 6.040 26.200 7.430 ;
        RECT 133.655 7.420 140.840 8.485 ;
        RECT 141.460 8.000 141.690 8.090 ;
        RECT 141.900 8.000 142.130 8.090 ;
        RECT 142.840 8.000 143.240 8.900 ;
        RECT 144.820 8.000 145.050 8.060 ;
        RECT 145.260 8.000 145.490 8.060 ;
        RECT 141.355 7.650 141.715 8.000 ;
        RECT 141.880 7.650 142.240 8.000 ;
        RECT 142.790 7.650 143.290 8.000 ;
        RECT 144.705 7.650 145.065 8.000 ;
        RECT 145.230 7.650 145.590 8.000 ;
        RECT 141.460 7.090 141.690 7.650 ;
        RECT 141.900 7.090 142.130 7.650 ;
        RECT 142.840 7.600 143.240 7.650 ;
        RECT 144.820 7.060 145.050 7.650 ;
        RECT 145.260 7.060 145.490 7.650 ;
        RECT 146.390 6.955 146.690 8.900 ;
        RECT 149.390 8.485 149.740 16.475 ;
        RECT 146.840 7.420 151.990 8.485 ;
        RECT 139.690 6.900 140.090 6.950 ;
        RECT 146.335 6.900 146.745 6.955 ;
        RECT 139.690 6.650 146.745 6.900 ;
        RECT 139.690 6.600 140.090 6.650 ;
        RECT 146.335 6.595 146.745 6.650 ;
      LAYER met2 ;
        RECT 22.630 223.785 22.910 224.155 ;
        RECT 4.230 222.425 4.510 222.795 ;
        RECT 7.910 222.425 8.190 222.795 ;
        RECT 11.590 222.425 11.870 222.795 ;
        RECT 16.190 222.425 16.470 222.795 ;
        RECT 18.950 222.425 19.230 222.795 ;
        RECT 22.700 222.600 22.840 223.785 ;
        RECT 78.760 223.640 79.020 223.960 ;
        RECT 79.210 223.785 79.490 224.155 ;
        RECT 85.190 223.785 85.470 224.155 ;
        RECT 40.860 222.855 42.400 223.225 ;
        RECT 48.390 223.105 48.670 223.475 ;
        RECT 4.240 222.280 4.500 222.425 ;
        RECT 7.920 222.280 8.180 222.425 ;
        RECT 11.600 222.280 11.860 222.425 ;
        RECT 16.200 222.280 16.460 222.425 ;
        RECT 18.960 222.280 19.220 222.425 ;
        RECT 22.640 222.280 22.900 222.600 ;
        RECT 26.310 222.425 26.590 222.795 ;
        RECT 29.990 222.425 30.270 222.795 ;
        RECT 26.320 222.280 26.580 222.425 ;
        RECT 30.000 222.280 30.260 222.425 ;
        RECT 48.460 222.260 48.600 223.105 ;
        RECT 69.560 222.280 69.820 222.600 ;
        RECT 70.470 222.425 70.750 222.795 ;
        RECT 70.480 222.280 70.740 222.425 ;
        RECT 78.300 222.280 78.560 222.600 ;
        RECT 48.400 221.940 48.660 222.260 ;
        RECT 63.120 221.705 63.380 222.025 ;
        RECT 66.800 221.940 67.060 222.260 ;
        RECT 62.660 220.920 62.920 221.240 ;
        RECT 1.030 220.135 2.570 220.505 ;
        RECT 21.425 220.135 22.965 220.505 ;
        RECT 60.295 220.135 61.835 220.505 ;
        RECT 56.680 218.540 56.940 218.860 ;
        RECT 57.600 218.540 57.860 218.860 ;
        RECT 56.220 218.200 56.480 218.520 ;
        RECT 40.860 217.415 42.400 217.785 ;
        RECT 1.030 214.695 2.570 215.065 ;
        RECT 21.425 214.695 22.965 215.065 ;
        RECT 55.760 214.120 56.020 214.440 ;
        RECT 55.820 213.955 55.960 214.120 ;
        RECT 55.750 213.585 56.030 213.955 ;
        RECT 40.860 211.975 42.400 212.345 ;
        RECT 11.600 211.060 11.860 211.380 ;
        RECT 19.420 211.060 19.680 211.380 ;
        RECT 55.820 211.235 55.960 213.585 ;
        RECT 9.300 210.040 9.560 210.360 ;
        RECT 1.030 209.255 2.570 209.625 ;
        RECT 9.360 208.320 9.500 210.040 ;
        RECT 9.300 208.000 9.560 208.320 ;
        RECT 11.660 207.980 11.800 211.060 ;
        RECT 17.120 210.720 17.380 211.040 ;
        RECT 11.600 207.660 11.860 207.980 ;
        RECT 15.280 207.320 15.540 207.640 ;
        RECT 15.340 205.940 15.480 207.320 ;
        RECT 17.180 206.280 17.320 210.720 ;
        RECT 19.480 207.980 19.620 211.060 ;
        RECT 55.750 210.865 56.030 211.235 ;
        RECT 56.280 210.555 56.420 218.200 ;
        RECT 56.740 216.140 56.880 218.540 ;
        RECT 56.680 215.820 56.940 216.140 ;
        RECT 56.740 211.380 56.880 215.820 ;
        RECT 57.660 211.720 57.800 218.540 ;
        RECT 58.980 215.480 59.240 215.800 ;
        RECT 57.600 211.400 57.860 211.720 ;
        RECT 56.680 211.060 56.940 211.380 ;
        RECT 20.800 210.040 21.060 210.360 ;
        RECT 56.210 210.185 56.490 210.555 ;
        RECT 59.040 210.110 59.180 215.480 ;
        RECT 60.295 214.695 61.835 215.065 ;
        RECT 62.200 214.120 62.460 214.440 ;
        RECT 59.890 212.905 60.170 213.275 ;
        RECT 59.960 210.360 60.100 212.905 ;
        RECT 60.820 212.760 61.080 213.080 ;
        RECT 61.740 212.760 62.000 213.080 ;
        RECT 60.880 211.380 61.020 212.760 ;
        RECT 61.800 211.720 61.940 212.760 ;
        RECT 62.260 211.915 62.400 214.120 ;
        RECT 62.720 213.420 62.860 220.920 ;
        RECT 63.180 216.140 63.320 221.705 ;
        RECT 66.860 221.580 67.000 221.940 ;
        RECT 67.720 221.830 67.980 221.920 ;
        RECT 69.100 221.830 69.360 222.000 ;
        RECT 67.720 221.690 69.360 221.830 ;
        RECT 67.720 221.600 67.980 221.690 ;
        RECT 69.100 221.680 69.360 221.690 ;
        RECT 66.340 221.260 66.600 221.580 ;
        RECT 66.800 221.260 67.060 221.580 ;
        RECT 65.880 220.920 66.140 221.240 ;
        RECT 65.940 218.520 66.080 220.920 ;
        RECT 65.880 218.200 66.140 218.520 ;
        RECT 65.940 216.820 66.080 218.200 ;
        RECT 65.880 216.500 66.140 216.820 ;
        RECT 66.400 216.480 66.540 221.260 ;
        RECT 65.420 216.160 65.680 216.480 ;
        RECT 66.340 216.160 66.600 216.480 ;
        RECT 63.120 215.820 63.380 216.140 ;
        RECT 63.180 214.100 63.320 215.820 ;
        RECT 65.480 214.440 65.620 216.160 ;
        RECT 67.780 216.140 67.920 221.600 ;
        RECT 69.100 220.920 69.360 221.240 ;
        RECT 67.720 215.820 67.980 216.140 ;
        RECT 65.420 214.120 65.680 214.440 ;
        RECT 63.120 213.780 63.380 214.100 ;
        RECT 66.800 213.780 67.060 214.100 ;
        RECT 62.660 213.100 62.920 213.420 ;
        RECT 61.740 211.400 62.000 211.720 ;
        RECT 62.190 211.545 62.470 211.915 ;
        RECT 60.820 211.060 61.080 211.380 ;
        RECT 20.860 207.980 21.000 210.040 ;
        RECT 58.980 209.790 59.240 210.110 ;
        RECT 59.900 210.040 60.160 210.360 ;
        RECT 21.425 209.255 22.965 209.625 ;
        RECT 60.295 209.255 61.835 209.625 ;
        RECT 59.430 208.825 59.710 209.195 ;
        RECT 26.320 208.000 26.580 208.320 ;
        RECT 19.420 207.660 19.680 207.980 ;
        RECT 20.800 207.660 21.060 207.980 ;
        RECT 17.120 205.960 17.380 206.280 ;
        RECT 10.670 205.570 10.950 205.795 ;
        RECT 15.280 205.620 15.540 205.940 ;
        RECT 19.480 205.600 19.620 207.660 ;
        RECT 26.380 207.640 26.520 208.000 ;
        RECT 58.520 207.660 58.780 207.980 ;
        RECT 26.320 207.320 26.580 207.640 ;
        RECT 11.600 205.570 11.860 205.600 ;
        RECT 10.670 205.310 11.860 205.570 ;
        RECT 11.600 205.280 11.860 205.310 ;
        RECT 19.420 205.280 19.680 205.600 ;
        RECT 21.710 205.570 21.990 205.795 ;
        RECT 26.380 205.600 26.520 207.320 ;
        RECT 40.860 206.535 42.400 206.905 ;
        RECT 58.580 206.475 58.720 207.660 ;
        RECT 59.500 207.640 59.640 208.825 ;
        RECT 61.740 208.680 62.000 209.000 ;
        RECT 61.800 207.980 61.940 208.680 ;
        RECT 61.740 207.660 62.000 207.980 ;
        RECT 59.440 207.320 59.700 207.640 ;
        RECT 32.760 205.960 33.020 206.280 ;
        RECT 40.120 205.960 40.380 206.280 ;
        RECT 58.510 206.105 58.790 206.475 ;
        RECT 58.980 205.960 59.240 206.280 ;
        RECT 32.820 205.795 32.960 205.960 ;
        RECT 40.180 205.795 40.320 205.960 ;
        RECT 59.040 205.795 59.180 205.960 ;
        RECT 61.800 205.940 61.940 207.660 ;
        RECT 22.640 205.570 22.900 205.600 ;
        RECT 21.710 205.310 22.900 205.570 ;
        RECT 22.640 205.280 22.900 205.310 ;
        RECT 26.320 205.280 26.580 205.600 ;
        RECT 32.750 205.425 33.030 205.795 ;
        RECT 33.680 205.280 33.940 205.600 ;
        RECT 40.110 205.425 40.390 205.795 ;
        RECT 58.970 205.425 59.250 205.795 ;
        RECT 61.740 205.620 62.000 205.940 ;
        RECT 1.030 203.815 2.570 204.185 ;
        RECT 21.425 203.815 22.965 204.185 ;
        RECT 33.740 202.200 33.880 205.280 ;
        RECT 60.295 203.815 61.835 204.185 ;
        RECT 62.260 202.540 62.400 211.545 ;
        RECT 63.180 210.990 63.320 213.780 ;
        RECT 64.960 213.275 65.220 213.420 ;
        RECT 64.950 212.905 65.230 213.275 ;
        RECT 65.420 213.100 65.680 213.420 ;
        RECT 64.500 211.400 64.760 211.720 ;
        RECT 63.180 210.850 63.780 210.990 ;
        RECT 63.120 210.380 63.380 210.700 ;
        RECT 63.640 210.530 63.780 210.850 ;
        RECT 62.650 207.465 62.930 207.835 ;
        RECT 62.720 205.600 62.860 207.465 ;
        RECT 63.180 205.795 63.320 210.380 ;
        RECT 63.580 210.210 63.840 210.530 ;
        RECT 64.560 208.055 64.700 211.400 ;
        RECT 64.960 210.040 65.220 210.360 ;
        RECT 65.020 208.055 65.160 210.040 ;
        RECT 65.480 208.515 65.620 213.100 ;
        RECT 66.860 211.040 67.000 213.780 ;
        RECT 67.260 213.175 67.520 213.495 ;
        RECT 67.320 211.720 67.460 213.175 ;
        RECT 67.780 213.080 67.920 215.820 ;
        RECT 67.720 212.760 67.980 213.080 ;
        RECT 67.780 211.720 67.920 212.760 ;
        RECT 69.160 211.720 69.300 220.920 ;
        RECT 67.260 211.400 67.520 211.720 ;
        RECT 67.720 211.400 67.980 211.720 ;
        RECT 69.100 211.400 69.360 211.720 ;
        RECT 66.800 210.720 67.060 211.040 ;
        RECT 69.100 210.040 69.360 210.360 ;
        RECT 65.410 208.145 65.690 208.515 ;
        RECT 66.330 208.145 66.610 208.515 ;
        RECT 68.180 208.230 68.440 208.320 ;
        RECT 64.500 207.735 64.760 208.055 ;
        RECT 64.960 207.835 65.220 208.055 ;
        RECT 65.420 208.000 65.680 208.145 ;
        RECT 64.950 207.465 65.230 207.835 ;
        RECT 66.400 207.640 66.540 208.145 ;
        RECT 68.180 208.090 68.840 208.230 ;
        RECT 69.160 208.120 69.300 210.040 ;
        RECT 68.180 208.000 68.440 208.090 ;
        RECT 68.700 207.640 68.840 208.090 ;
        RECT 69.100 207.800 69.360 208.120 ;
        RECT 66.340 207.320 66.600 207.640 ;
        RECT 68.180 207.320 68.440 207.640 ;
        RECT 68.640 207.320 68.900 207.640 ;
        RECT 62.660 205.280 62.920 205.600 ;
        RECT 63.110 205.425 63.390 205.795 ;
        RECT 68.240 205.700 68.380 207.320 ;
        RECT 69.160 205.940 69.300 207.800 ;
        RECT 63.120 205.280 63.380 205.425 ;
        RECT 68.180 205.380 68.440 205.700 ;
        RECT 69.100 205.620 69.360 205.940 ;
        RECT 69.620 205.260 69.760 222.280 ;
        RECT 71.860 221.940 72.120 222.260 ;
        RECT 71.400 221.600 71.660 221.920 ;
        RECT 70.010 219.025 70.290 219.395 ;
        RECT 70.020 218.880 70.280 219.025 ;
        RECT 70.080 218.520 70.220 218.880 ;
        RECT 70.940 218.540 71.200 218.860 ;
        RECT 70.020 218.200 70.280 218.520 ;
        RECT 71.000 217.160 71.140 218.540 ;
        RECT 70.940 216.840 71.200 217.160 ;
        RECT 70.930 216.305 71.210 216.675 ;
        RECT 71.000 213.080 71.140 216.305 ;
        RECT 70.940 212.760 71.200 213.080 ;
        RECT 71.460 212.390 71.600 221.600 ;
        RECT 71.920 218.935 72.060 221.940 ;
        RECT 73.690 221.745 73.970 222.115 ;
        RECT 71.860 218.615 72.120 218.935 ;
        RECT 73.760 218.520 73.900 221.745 ;
        RECT 77.840 221.720 78.100 222.040 ;
        RECT 74.620 221.260 74.880 221.580 ;
        RECT 77.380 221.260 77.640 221.580 ;
        RECT 72.320 218.200 72.580 218.520 ;
        RECT 73.700 218.200 73.960 218.520 ;
        RECT 71.860 216.160 72.120 216.480 ;
        RECT 71.920 213.275 72.060 216.160 ;
        RECT 71.850 212.905 72.130 213.275 ;
        RECT 71.000 212.250 71.600 212.390 ;
        RECT 70.020 211.060 70.280 211.380 ;
        RECT 70.080 207.980 70.220 211.060 ;
        RECT 71.000 211.040 71.140 212.250 ;
        RECT 71.400 211.400 71.660 211.720 ;
        RECT 70.940 210.720 71.200 211.040 ;
        RECT 71.000 207.980 71.140 210.720 ;
        RECT 71.460 210.110 71.600 211.400 ;
        RECT 71.920 211.040 72.060 212.905 ;
        RECT 72.380 211.720 72.520 218.200 ;
        RECT 74.680 216.675 74.820 221.260 ;
        RECT 77.440 218.860 77.580 221.260 ;
        RECT 77.900 218.860 78.040 221.720 ;
        RECT 78.360 221.490 78.500 222.280 ;
        RECT 78.820 222.090 78.960 223.640 ;
        RECT 78.760 221.770 79.020 222.090 ;
        RECT 78.360 221.350 78.960 221.490 ;
        RECT 75.600 218.705 76.660 218.845 ;
        RECT 74.610 216.305 74.890 216.675 ;
        RECT 74.620 216.160 74.880 216.305 ;
        RECT 74.680 213.760 74.820 216.160 ;
        RECT 74.620 213.440 74.880 213.760 ;
        RECT 75.080 213.440 75.340 213.760 ;
        RECT 72.320 211.400 72.580 211.720 ;
        RECT 71.860 210.720 72.120 211.040 ;
        RECT 71.400 209.790 71.660 210.110 ;
        RECT 74.160 210.040 74.420 210.360 ;
        RECT 70.020 207.835 70.280 207.980 ;
        RECT 70.010 207.465 70.290 207.835 ;
        RECT 70.940 207.660 71.200 207.980 ;
        RECT 71.460 205.940 71.600 209.790 ;
        RECT 72.780 208.680 73.040 209.000 ;
        RECT 71.400 205.795 71.660 205.940 ;
        RECT 71.390 205.425 71.670 205.795 ;
        RECT 72.840 205.705 72.980 208.680 ;
        RECT 74.220 206.280 74.360 210.040 ;
        RECT 75.140 208.660 75.280 213.440 ;
        RECT 75.600 211.040 75.740 218.705 ;
        RECT 76.520 218.520 76.660 218.705 ;
        RECT 76.920 218.540 77.180 218.860 ;
        RECT 77.380 218.540 77.640 218.860 ;
        RECT 77.840 218.540 78.100 218.860 ;
        RECT 76.000 218.200 76.260 218.520 ;
        RECT 76.460 218.200 76.720 218.520 ;
        RECT 76.060 215.800 76.200 218.200 ;
        RECT 76.980 216.480 77.120 218.540 ;
        RECT 76.920 216.160 77.180 216.480 ;
        RECT 76.460 215.820 76.720 216.140 ;
        RECT 76.000 215.480 76.260 215.800 ;
        RECT 76.060 213.420 76.200 215.480 ;
        RECT 76.520 213.420 76.660 215.820 ;
        RECT 76.920 213.780 77.180 214.100 ;
        RECT 76.000 213.100 76.260 213.420 ;
        RECT 76.460 213.100 76.720 213.420 ;
        RECT 76.980 213.080 77.120 213.780 ;
        RECT 78.300 213.100 78.560 213.420 ;
        RECT 78.820 213.275 78.960 221.350 ;
        RECT 76.920 212.760 77.180 213.080 ;
        RECT 76.980 211.145 77.120 212.760 ;
        RECT 78.360 212.480 78.500 213.100 ;
        RECT 78.750 212.905 79.030 213.275 ;
        RECT 79.280 212.480 79.420 223.785 ;
        RECT 79.730 222.855 81.270 223.225 ;
        RECT 85.260 222.260 85.400 223.785 ;
        RECT 116.480 223.640 116.740 223.960 ;
        RECT 117.400 223.640 117.660 223.960 ;
        RECT 126.130 223.785 126.410 224.155 ;
        RECT 89.340 222.280 89.600 222.600 ;
        RECT 95.780 222.510 96.040 222.600 ;
        RECT 94.920 222.370 96.040 222.510 ;
        RECT 81.520 221.705 81.780 222.025 ;
        RECT 84.280 221.705 84.540 222.025 ;
        RECT 85.200 221.940 85.460 222.260 ;
        RECT 79.730 217.415 81.270 217.785 ;
        RECT 81.580 215.880 81.720 221.705 ;
        RECT 81.980 220.920 82.240 221.240 ;
        RECT 82.900 220.920 83.160 221.240 ;
        RECT 82.040 216.820 82.180 220.920 ;
        RECT 82.960 218.860 83.100 220.920 ;
        RECT 82.900 218.540 83.160 218.860 ;
        RECT 81.980 216.500 82.240 216.820 ;
        RECT 80.660 215.800 81.720 215.880 ;
        RECT 80.600 215.740 81.720 215.800 ;
        RECT 80.600 215.480 80.860 215.740 ;
        RECT 81.580 213.495 81.720 215.740 ;
        RECT 81.520 213.175 81.780 213.495 ;
        RECT 78.360 212.340 79.420 212.480 ;
        RECT 79.730 211.975 81.270 212.345 ;
        RECT 81.980 211.400 82.240 211.720 ;
        RECT 75.540 210.950 75.800 211.040 ;
        RECT 75.540 210.810 76.200 210.950 ;
        RECT 76.920 210.825 77.180 211.145 ;
        RECT 78.300 210.825 78.560 211.145 ;
        RECT 75.540 210.720 75.800 210.810 ;
        RECT 75.530 209.505 75.810 209.875 ;
        RECT 75.080 208.340 75.340 208.660 ;
        RECT 75.600 208.065 75.740 209.505 ;
        RECT 76.060 209.195 76.200 210.810 ;
        RECT 77.380 210.380 77.640 210.700 ;
        RECT 77.840 210.555 78.100 210.700 ;
        RECT 75.990 208.825 76.270 209.195 ;
        RECT 75.540 207.745 75.800 208.065 ;
        RECT 76.920 208.000 77.180 208.320 ;
        RECT 74.160 205.960 74.420 206.280 ;
        RECT 71.860 205.280 72.120 205.600 ;
        RECT 72.780 205.385 73.040 205.705 ;
        RECT 69.560 204.940 69.820 205.260 ;
        RECT 62.200 202.220 62.460 202.540 ;
        RECT 33.680 201.880 33.940 202.200 ;
        RECT 64.040 201.880 64.300 202.200 ;
        RECT 40.860 201.095 42.400 201.465 ;
        RECT 64.100 200.355 64.240 201.880 ;
        RECT 71.920 201.035 72.060 205.280 ;
        RECT 76.000 204.940 76.260 205.260 ;
        RECT 76.060 202.615 76.200 204.940 ;
        RECT 76.980 203.220 77.120 208.000 ;
        RECT 77.440 205.600 77.580 210.380 ;
        RECT 77.830 210.185 78.110 210.555 ;
        RECT 77.840 205.960 78.100 206.280 ;
        RECT 77.900 205.795 78.040 205.960 ;
        RECT 77.380 205.280 77.640 205.600 ;
        RECT 77.830 205.425 78.110 205.795 ;
        RECT 76.920 202.900 77.180 203.220 ;
        RECT 78.360 202.615 78.500 210.825 ;
        RECT 81.050 210.185 81.330 210.555 ;
        RECT 81.120 208.320 81.260 210.185 ;
        RECT 81.520 208.910 81.780 209.000 ;
        RECT 82.040 208.910 82.180 211.400 ;
        RECT 84.340 210.700 84.480 221.705 ;
        RECT 86.120 221.600 86.380 221.920 ;
        RECT 87.030 221.745 87.310 222.115 ;
        RECT 86.180 219.880 86.320 221.600 ;
        RECT 86.120 219.790 86.380 219.880 ;
        RECT 85.720 219.650 86.380 219.790 ;
        RECT 85.720 216.675 85.860 219.650 ;
        RECT 86.120 219.560 86.380 219.650 ;
        RECT 87.100 219.200 87.240 221.745 ;
        RECT 87.040 218.880 87.300 219.200 ;
        RECT 89.400 218.935 89.540 222.280 ;
        RECT 94.920 221.920 95.060 222.370 ;
        RECT 95.780 222.280 96.040 222.370 ;
        RECT 98.080 222.280 98.340 222.600 ;
        RECT 94.860 221.600 95.120 221.920 ;
        RECT 95.320 221.640 95.580 221.960 ;
        RECT 96.240 221.640 96.500 221.960 ;
        RECT 95.380 219.540 95.520 221.640 ;
        RECT 95.320 219.220 95.580 219.540 ;
        RECT 87.960 218.615 88.220 218.935 ;
        RECT 89.340 218.615 89.600 218.935 ;
        RECT 89.800 218.880 90.060 219.200 ;
        RECT 85.650 216.305 85.930 216.675 ;
        RECT 85.200 215.710 85.460 215.800 ;
        RECT 84.800 215.570 85.460 215.710 ;
        RECT 84.800 213.760 84.940 215.570 ;
        RECT 85.200 215.480 85.460 215.570 ;
        RECT 84.740 213.440 85.000 213.760 ;
        RECT 85.190 213.585 85.470 213.955 ;
        RECT 84.800 211.120 84.940 213.440 ;
        RECT 84.740 210.800 85.000 211.120 ;
        RECT 82.900 210.380 83.160 210.700 ;
        RECT 84.280 210.380 84.540 210.700 ;
        RECT 81.520 208.770 82.180 208.910 ;
        RECT 82.430 208.825 82.710 209.195 ;
        RECT 81.520 208.680 81.780 208.770 ;
        RECT 81.060 208.000 81.320 208.320 ;
        RECT 78.760 207.320 79.020 207.640 ;
        RECT 79.220 207.320 79.480 207.640 ;
        RECT 76.000 202.295 76.260 202.615 ;
        RECT 78.300 202.295 78.560 202.615 ;
        RECT 78.820 202.540 78.960 207.320 ;
        RECT 79.280 205.940 79.420 207.320 ;
        RECT 79.730 206.535 81.270 206.905 ;
        RECT 79.220 205.620 79.480 205.940 ;
        RECT 80.590 205.425 80.870 205.795 ;
        RECT 82.500 205.705 82.640 208.825 ;
        RECT 82.960 208.660 83.100 210.380 ;
        RECT 84.340 209.080 84.480 210.380 ;
        RECT 83.420 208.940 84.480 209.080 ;
        RECT 84.800 209.000 84.940 210.800 ;
        RECT 82.900 208.340 83.160 208.660 ;
        RECT 83.420 206.280 83.560 208.940 ;
        RECT 84.740 208.680 85.000 209.000 ;
        RECT 84.280 208.000 84.540 208.320 ;
        RECT 84.740 208.000 85.000 208.320 ;
        RECT 84.340 207.155 84.480 208.000 ;
        RECT 84.270 206.785 84.550 207.155 ;
        RECT 83.360 205.960 83.620 206.280 ;
        RECT 80.660 205.260 80.800 205.425 ;
        RECT 82.440 205.385 82.700 205.705 ;
        RECT 80.600 204.940 80.860 205.260 ;
        RECT 84.800 203.220 84.940 208.000 ;
        RECT 85.260 207.890 85.400 213.585 ;
        RECT 85.720 211.040 85.860 216.305 ;
        RECT 86.580 215.820 86.840 216.140 ;
        RECT 86.640 213.080 86.780 215.820 ;
        RECT 86.580 212.760 86.840 213.080 ;
        RECT 85.660 210.720 85.920 211.040 ;
        RECT 86.110 210.865 86.390 211.235 ;
        RECT 86.640 211.160 86.780 212.760 ;
        RECT 85.720 210.555 85.860 210.720 ;
        RECT 85.650 210.185 85.930 210.555 ;
        RECT 86.180 209.000 86.320 210.865 ;
        RECT 86.580 210.840 86.840 211.160 ;
        RECT 87.040 211.060 87.300 211.380 ;
        RECT 86.120 208.680 86.380 209.000 ;
        RECT 85.660 207.890 85.920 207.980 ;
        RECT 85.260 207.750 85.920 207.890 ;
        RECT 85.660 207.660 85.920 207.750 ;
        RECT 86.120 207.320 86.380 207.640 ;
        RECT 86.180 205.705 86.320 207.320 ;
        RECT 86.640 207.155 86.780 210.840 ;
        RECT 87.100 209.875 87.240 211.060 ;
        RECT 87.030 209.505 87.310 209.875 ;
        RECT 88.020 207.980 88.160 218.615 ;
        RECT 89.860 216.140 90.000 218.880 ;
        RECT 93.940 218.200 94.200 218.520 ;
        RECT 94.000 216.820 94.140 218.200 ;
        RECT 96.300 217.160 96.440 221.640 ;
        RECT 96.700 220.920 96.960 221.240 ;
        RECT 96.760 217.160 96.900 220.920 ;
        RECT 98.140 218.860 98.280 222.280 ;
        RECT 109.120 221.940 109.380 222.260 ;
        RECT 108.660 221.260 108.920 221.580 ;
        RECT 108.200 220.920 108.460 221.240 ;
        RECT 99.165 220.135 100.705 220.505 ;
        RECT 99.460 219.220 99.720 219.540 ;
        RECT 98.540 218.880 98.800 219.200 ;
        RECT 98.080 218.540 98.340 218.860 ;
        RECT 96.240 216.840 96.500 217.160 ;
        RECT 96.700 216.840 96.960 217.160 ;
        RECT 93.940 216.500 94.200 216.820 ;
        RECT 96.300 216.480 96.440 216.840 ;
        RECT 98.080 216.670 98.340 216.990 ;
        RECT 96.240 216.160 96.500 216.480 ;
        RECT 89.800 215.820 90.060 216.140 ;
        RECT 98.140 213.760 98.280 216.670 ;
        RECT 98.080 213.440 98.340 213.760 ;
        RECT 91.170 212.905 91.450 213.275 ;
        RECT 91.180 212.760 91.440 212.905 ;
        RECT 90.260 210.380 90.520 210.700 ;
        RECT 96.240 210.380 96.500 210.700 ;
        RECT 97.160 210.555 97.420 210.700 ;
        RECT 90.320 208.660 90.460 210.380 ;
        RECT 90.260 208.340 90.520 208.660 ;
        RECT 96.300 208.320 96.440 210.380 ;
        RECT 97.150 210.185 97.430 210.555 ;
        RECT 98.600 208.320 98.740 218.880 ;
        RECT 99.520 218.860 99.660 219.220 ;
        RECT 108.260 219.200 108.400 220.920 ;
        RECT 108.720 220.075 108.860 221.260 ;
        RECT 108.650 219.705 108.930 220.075 ;
        RECT 108.200 218.880 108.460 219.200 ;
        RECT 99.460 218.540 99.720 218.860 ;
        RECT 99.520 215.995 99.660 218.540 ;
        RECT 107.280 216.160 107.540 216.480 ;
        RECT 99.450 215.625 99.730 215.995 ;
        RECT 99.165 214.695 100.705 215.065 ;
        RECT 107.340 214.440 107.480 216.160 ;
        RECT 107.280 214.120 107.540 214.440 ;
        RECT 104.580 213.760 105.640 213.840 ;
        RECT 104.520 213.700 105.700 213.760 ;
        RECT 104.520 213.440 104.780 213.700 ;
        RECT 105.440 213.440 105.700 213.700 ;
        RECT 99.460 212.760 99.720 213.080 ;
        RECT 104.060 212.760 104.320 213.080 ;
        RECT 105.900 212.990 106.160 213.080 ;
        RECT 107.280 212.990 107.540 213.080 ;
        RECT 105.900 212.850 107.540 212.990 ;
        RECT 105.900 212.760 106.160 212.850 ;
        RECT 107.280 212.760 107.540 212.850 ;
        RECT 99.000 211.235 99.260 211.380 ;
        RECT 98.990 210.865 99.270 211.235 ;
        RECT 99.520 211.040 99.660 212.760 ;
        RECT 101.300 211.235 101.560 211.380 ;
        RECT 99.460 210.720 99.720 211.040 ;
        RECT 101.290 210.865 101.570 211.235 ;
        RECT 101.760 211.060 102.020 211.380 ;
        RECT 100.380 210.270 100.640 210.360 ;
        RECT 100.380 210.130 101.040 210.270 ;
        RECT 100.380 210.040 100.640 210.130 ;
        RECT 99.165 209.255 100.705 209.625 ;
        RECT 96.240 208.000 96.500 208.320 ;
        RECT 98.540 208.000 98.800 208.320 ;
        RECT 87.490 207.465 87.770 207.835 ;
        RECT 87.960 207.660 88.220 207.980 ;
        RECT 88.420 207.660 88.680 207.980 ;
        RECT 86.570 206.785 86.850 207.155 ;
        RECT 87.560 205.940 87.700 207.465 ;
        RECT 86.120 205.385 86.380 205.705 ;
        RECT 87.500 205.620 87.760 205.940 ;
        RECT 88.480 205.795 88.620 207.660 ;
        RECT 100.900 207.640 101.040 210.130 ;
        RECT 101.820 208.515 101.960 211.060 ;
        RECT 104.120 210.700 104.260 212.760 ;
        RECT 104.970 210.865 105.250 211.235 ;
        RECT 107.340 211.210 107.480 212.760 ;
        RECT 108.260 211.380 108.400 218.880 ;
        RECT 109.180 214.440 109.320 221.940 ;
        RECT 109.580 221.830 109.840 221.920 ;
        RECT 110.500 221.830 110.760 221.920 ;
        RECT 109.580 221.690 110.760 221.830 ;
        RECT 109.580 221.600 109.840 221.690 ;
        RECT 110.500 221.600 110.760 221.690 ;
        RECT 115.100 221.600 115.360 221.920 ;
        RECT 116.020 221.600 116.280 221.920 ;
        RECT 109.640 219.540 109.780 221.600 ;
        RECT 110.040 220.920 110.300 221.240 ;
        RECT 110.500 220.920 110.760 221.240 ;
        RECT 110.100 219.880 110.240 220.920 ;
        RECT 110.040 219.560 110.300 219.880 ;
        RECT 109.580 219.220 109.840 219.540 ;
        RECT 109.120 214.120 109.380 214.440 ;
        RECT 109.120 213.440 109.380 213.760 ;
        RECT 107.280 210.890 107.540 211.210 ;
        RECT 108.200 211.060 108.460 211.380 ;
        RECT 104.060 210.555 104.320 210.700 ;
        RECT 103.600 210.040 103.860 210.360 ;
        RECT 104.050 210.185 104.330 210.555 ;
        RECT 104.520 210.040 104.780 210.360 ;
        RECT 101.750 208.145 102.030 208.515 ;
        RECT 88.880 207.320 89.140 207.640 ;
        RECT 96.240 207.320 96.500 207.640 ;
        RECT 98.080 207.320 98.340 207.640 ;
        RECT 100.840 207.320 101.100 207.640 ;
        RECT 88.410 205.425 88.690 205.795 ;
        RECT 88.940 205.600 89.080 207.320 ;
        RECT 89.800 205.960 90.060 206.280 ;
        RECT 89.860 205.795 90.000 205.960 ;
        RECT 96.300 205.940 96.440 207.320 ;
        RECT 88.880 205.280 89.140 205.600 ;
        RECT 89.790 205.425 90.070 205.795 ;
        RECT 96.240 205.620 96.500 205.940 ;
        RECT 98.140 205.600 98.280 207.320 ;
        RECT 103.140 205.960 103.400 206.280 ;
        RECT 103.200 205.795 103.340 205.960 ;
        RECT 103.660 205.940 103.800 210.040 ;
        RECT 98.080 205.280 98.340 205.600 ;
        RECT 103.130 205.425 103.410 205.795 ;
        RECT 103.600 205.620 103.860 205.940 ;
        RECT 104.580 205.600 104.720 210.040 ;
        RECT 105.040 209.000 105.180 210.865 ;
        RECT 109.180 210.700 109.320 213.440 ;
        RECT 109.580 211.120 109.840 211.210 ;
        RECT 110.560 211.120 110.700 220.920 ;
        RECT 114.640 218.880 114.900 219.200 ;
        RECT 113.260 218.540 113.520 218.860 ;
        RECT 113.320 217.160 113.460 218.540 ;
        RECT 114.700 218.520 114.840 218.880 ;
        RECT 115.160 218.520 115.300 221.600 ;
        RECT 116.080 219.540 116.220 221.600 ;
        RECT 116.020 219.220 116.280 219.540 ;
        RECT 116.080 218.520 116.220 219.220 ;
        RECT 114.640 218.200 114.900 218.520 ;
        RECT 115.100 218.200 115.360 218.520 ;
        RECT 116.020 218.200 116.280 218.520 ;
        RECT 114.700 217.160 114.840 218.200 ;
        RECT 113.260 216.840 113.520 217.160 ;
        RECT 114.640 216.840 114.900 217.160 ;
        RECT 112.330 215.625 112.610 215.995 ;
        RECT 111.880 213.100 112.140 213.420 ;
        RECT 109.580 210.980 110.700 211.120 ;
        RECT 111.420 211.060 111.680 211.380 ;
        RECT 111.940 211.120 112.080 213.100 ;
        RECT 112.400 211.120 112.540 215.625 ;
        RECT 112.800 215.480 113.060 215.800 ;
        RECT 112.860 213.760 113.000 215.480 ;
        RECT 112.800 213.440 113.060 213.760 ;
        RECT 113.320 211.235 113.460 216.840 ;
        RECT 115.160 213.080 115.300 218.200 ;
        RECT 116.080 216.820 116.220 218.200 ;
        RECT 116.020 216.500 116.280 216.820 ;
        RECT 116.080 213.420 116.220 216.500 ;
        RECT 116.020 213.100 116.280 213.420 ;
        RECT 113.720 212.760 113.980 213.080 ;
        RECT 115.100 212.760 115.360 213.080 ;
        RECT 113.780 211.720 113.920 212.760 ;
        RECT 113.720 211.400 113.980 211.720 ;
        RECT 109.580 210.890 109.840 210.980 ;
        RECT 105.440 210.380 105.700 210.700 ;
        RECT 109.120 210.380 109.380 210.700 ;
        RECT 104.980 208.680 105.240 209.000 ;
        RECT 105.500 208.660 105.640 210.380 ;
        RECT 106.820 210.040 107.080 210.360 ;
        RECT 105.440 208.340 105.700 208.660 ;
        RECT 106.880 207.980 107.020 210.040 ;
        RECT 111.480 208.660 111.620 211.060 ;
        RECT 111.880 210.800 112.140 211.120 ;
        RECT 112.340 210.800 112.600 211.120 ;
        RECT 113.250 210.865 113.530 211.235 ;
        RECT 116.080 211.040 116.220 213.100 ;
        RECT 116.540 211.720 116.680 223.640 ;
        RECT 116.940 218.540 117.200 218.860 ;
        RECT 117.000 217.160 117.140 218.540 ;
        RECT 116.940 216.840 117.200 217.160 ;
        RECT 117.460 213.760 117.600 223.640 ;
        RECT 118.600 222.855 120.140 223.225 ;
        RECT 126.200 221.920 126.340 223.785 ;
        RECT 151.900 223.640 152.160 223.960 ;
        RECT 127.510 223.105 127.790 223.475 ;
        RECT 133.950 223.105 134.230 223.475 ;
        RECT 143.150 223.105 143.430 223.475 ;
        RECT 127.580 221.920 127.720 223.105 ;
        RECT 132.580 221.940 132.840 222.260 ;
        RECT 126.140 221.600 126.400 221.920 ;
        RECT 127.520 221.600 127.780 221.920 ;
        RECT 120.620 221.260 120.880 221.580 ;
        RECT 131.200 221.260 131.460 221.580 ;
        RECT 118.310 219.705 118.590 220.075 ;
        RECT 118.320 219.560 118.580 219.705 ;
        RECT 117.860 218.200 118.120 218.520 ;
        RECT 117.920 216.480 118.060 218.200 ;
        RECT 118.600 217.415 120.140 217.785 ;
        RECT 119.700 216.500 119.960 216.820 ;
        RECT 117.860 216.160 118.120 216.480 ;
        RECT 117.400 213.440 117.660 213.760 ;
        RECT 119.760 213.420 119.900 216.500 ;
        RECT 120.680 214.100 120.820 221.260 ;
        RECT 122.920 218.540 123.180 218.860 ;
        RECT 122.000 218.200 122.260 218.520 ;
        RECT 120.620 213.780 120.880 214.100 ;
        RECT 122.060 213.760 122.200 218.200 ;
        RECT 122.980 216.730 123.120 218.540 ;
        RECT 127.520 218.200 127.780 218.520 ;
        RECT 127.580 216.820 127.720 218.200 ;
        RECT 123.380 216.730 123.640 216.820 ;
        RECT 122.980 216.590 123.640 216.730 ;
        RECT 123.380 216.500 123.640 216.590 ;
        RECT 126.140 216.200 126.400 216.520 ;
        RECT 127.520 216.500 127.780 216.820 ;
        RECT 125.220 216.050 125.480 216.140 ;
        RECT 123.440 215.910 125.480 216.050 ;
        RECT 126.200 215.995 126.340 216.200 ;
        RECT 131.260 216.140 131.400 221.260 ;
        RECT 132.640 216.480 132.780 221.940 ;
        RECT 134.020 221.920 134.160 223.105 ;
        RECT 143.220 221.920 143.360 223.105 ;
        RECT 151.960 222.680 152.100 223.640 ;
        RECT 157.470 222.855 159.010 223.225 ;
        RECT 151.960 222.540 153.020 222.680 ;
        RECT 133.960 221.600 134.220 221.920 ;
        RECT 139.940 221.600 140.200 221.920 ;
        RECT 143.160 221.600 143.420 221.920 ;
        RECT 137.640 221.260 137.900 221.580 ;
        RECT 133.040 220.920 133.300 221.240 ;
        RECT 135.340 220.920 135.600 221.240 ;
        RECT 133.100 217.160 133.240 220.920 ;
        RECT 134.420 218.540 134.680 218.860 ;
        RECT 134.480 217.160 134.620 218.540 ;
        RECT 133.040 216.840 133.300 217.160 ;
        RECT 134.420 216.840 134.680 217.160 ;
        RECT 135.400 216.480 135.540 220.920 ;
        RECT 137.700 219.880 137.840 221.260 ;
        RECT 138.035 220.135 139.575 220.505 ;
        RECT 137.640 219.560 137.900 219.880 ;
        RECT 140.000 218.520 140.140 221.600 ;
        RECT 145.920 221.260 146.180 221.580 ;
        RECT 140.390 220.385 140.670 220.755 ;
        RECT 140.460 219.880 140.600 220.385 ;
        RECT 140.400 219.560 140.660 219.880 ;
        RECT 144.540 219.560 144.800 219.880 ;
        RECT 144.070 219.025 144.350 219.395 ;
        RECT 139.940 218.200 140.200 218.520 ;
        RECT 141.780 218.200 142.040 218.520 ;
        RECT 143.160 218.200 143.420 218.520 ;
        RECT 140.000 216.820 140.140 218.200 ;
        RECT 141.840 217.160 141.980 218.200 ;
        RECT 141.780 216.840 142.040 217.160 ;
        RECT 139.940 216.500 140.200 216.820 ;
        RECT 132.580 216.160 132.840 216.480 ;
        RECT 135.340 216.160 135.600 216.480 ;
        RECT 130.280 215.995 130.540 216.140 ;
        RECT 122.000 213.670 122.260 213.760 ;
        RECT 121.140 213.530 122.260 213.670 ;
        RECT 119.700 213.100 119.960 213.420 ;
        RECT 117.400 212.760 117.660 213.080 ;
        RECT 116.480 211.400 116.740 211.720 ;
        RECT 113.320 210.700 113.460 210.865 ;
        RECT 116.020 210.720 116.280 211.040 ;
        RECT 113.260 210.380 113.520 210.700 ;
        RECT 112.340 210.040 112.600 210.360 ;
        RECT 111.420 208.340 111.680 208.660 ;
        RECT 112.400 208.055 112.540 210.040 ;
        RECT 106.820 207.660 107.080 207.980 ;
        RECT 107.280 207.835 107.540 207.980 ;
        RECT 107.270 207.465 107.550 207.835 ;
        RECT 112.340 207.735 112.600 208.055 ;
        RECT 117.460 207.980 117.600 212.760 ;
        RECT 118.600 211.975 120.140 212.345 ;
        RECT 121.140 211.040 121.280 213.530 ;
        RECT 122.000 213.440 122.260 213.530 ;
        RECT 122.460 213.100 122.720 213.420 ;
        RECT 122.520 212.390 122.660 213.100 ;
        RECT 123.440 212.390 123.580 215.910 ;
        RECT 125.220 215.820 125.480 215.910 ;
        RECT 126.130 215.625 126.410 215.995 ;
        RECT 130.270 215.625 130.550 215.995 ;
        RECT 131.200 215.820 131.460 216.140 ;
        RECT 137.180 215.820 137.440 216.140 ;
        RECT 130.340 213.420 130.480 215.625 ;
        RECT 132.120 215.480 132.380 215.800 ;
        RECT 132.180 214.440 132.320 215.480 ;
        RECT 132.120 214.120 132.380 214.440 ;
        RECT 137.240 213.760 137.380 215.820 ;
        RECT 138.035 214.695 139.575 215.065 ;
        RECT 143.220 214.440 143.360 218.200 ;
        RECT 143.160 214.120 143.420 214.440 ;
        RECT 137.180 213.440 137.440 213.760 ;
        RECT 144.140 213.420 144.280 219.025 ;
        RECT 144.600 216.480 144.740 219.560 ;
        RECT 145.000 218.540 145.260 218.860 ;
        RECT 144.540 216.160 144.800 216.480 ;
        RECT 145.060 216.140 145.200 218.540 ;
        RECT 145.000 215.820 145.260 216.140 ;
        RECT 145.980 214.440 146.120 221.260 ;
        RECT 147.300 220.920 147.560 221.240 ;
        RECT 146.380 218.540 146.640 218.860 ;
        RECT 146.440 214.440 146.580 218.540 ;
        RECT 146.840 218.200 147.100 218.520 ;
        RECT 146.900 216.480 147.040 218.200 ;
        RECT 146.840 216.160 147.100 216.480 ;
        RECT 145.920 214.120 146.180 214.440 ;
        RECT 146.380 214.120 146.640 214.440 ;
        RECT 147.360 213.420 147.500 220.920 ;
        RECT 147.750 220.385 148.030 220.755 ;
        RECT 147.820 217.160 147.960 220.385 ;
        RECT 151.960 219.880 152.100 222.540 ;
        RECT 152.880 221.920 153.020 222.540 ;
        RECT 155.580 222.280 155.840 222.600 ;
        RECT 152.360 221.600 152.620 221.920 ;
        RECT 152.820 221.600 153.080 221.920 ;
        RECT 152.420 219.880 152.560 221.600 ;
        RECT 154.200 221.260 154.460 221.580 ;
        RECT 152.820 220.920 153.080 221.240 ;
        RECT 151.900 219.560 152.160 219.880 ;
        RECT 152.360 219.560 152.620 219.880 ;
        RECT 147.760 216.840 148.020 217.160 ;
        RECT 152.360 216.500 152.620 216.820 ;
        RECT 152.420 214.440 152.560 216.500 ;
        RECT 152.360 214.120 152.620 214.440 ;
        RECT 152.880 213.420 153.020 220.920 ;
        RECT 154.260 217.160 154.400 221.260 ;
        RECT 154.650 219.705 154.930 220.075 ;
        RECT 154.200 216.840 154.460 217.160 ;
        RECT 154.720 214.100 154.860 219.705 ;
        RECT 155.640 219.200 155.780 222.280 ;
        RECT 155.580 218.880 155.840 219.200 ;
        RECT 155.640 215.800 155.780 218.880 ;
        RECT 157.470 217.415 159.010 217.785 ;
        RECT 155.580 215.480 155.840 215.800 ;
        RECT 154.660 213.780 154.920 214.100 ;
        RECT 130.280 213.100 130.540 213.420 ;
        RECT 133.960 213.100 134.220 213.420 ;
        RECT 144.080 213.100 144.340 213.420 ;
        RECT 147.300 213.100 147.560 213.420 ;
        RECT 152.820 213.100 153.080 213.420 ;
        RECT 129.360 212.760 129.620 213.080 ;
        RECT 121.600 212.250 122.660 212.390 ;
        RECT 122.980 212.250 123.580 212.390 ;
        RECT 121.600 211.720 121.740 212.250 ;
        RECT 121.540 211.400 121.800 211.720 ;
        RECT 122.980 211.380 123.120 212.250 ;
        RECT 129.420 211.720 129.560 212.760 ;
        RECT 127.060 211.400 127.320 211.720 ;
        RECT 129.360 211.400 129.620 211.720 ;
        RECT 122.920 211.060 123.180 211.380 ;
        RECT 121.080 210.720 121.340 211.040 ;
        RECT 127.120 208.120 127.260 211.400 ;
        RECT 128.440 210.040 128.700 210.360 ;
        RECT 128.500 209.050 128.640 210.040 ;
        RECT 128.440 208.730 128.700 209.050 ;
        RECT 134.020 209.000 134.160 213.100 ;
        RECT 157.470 211.975 159.010 212.345 ;
        RECT 138.035 209.255 139.575 209.625 ;
        RECT 133.960 208.680 134.220 209.000 ;
        RECT 153.730 208.825 154.010 209.195 ;
        RECT 117.400 207.660 117.660 207.980 ;
        RECT 127.060 207.800 127.320 208.120 ;
        RECT 109.120 207.320 109.380 207.640 ;
        RECT 109.180 205.940 109.320 207.320 ;
        RECT 118.600 206.535 120.140 206.905 ;
        RECT 109.120 205.620 109.380 205.940 ;
        RECT 114.180 205.795 114.440 205.940 ;
        RECT 150.980 205.795 151.240 205.940 ;
        RECT 104.520 205.280 104.780 205.600 ;
        RECT 114.170 205.425 114.450 205.795 ;
        RECT 117.850 205.425 118.130 205.795 ;
        RECT 128.890 205.425 129.170 205.795 ;
        RECT 150.970 205.425 151.250 205.795 ;
        RECT 153.800 205.685 153.940 208.825 ;
        RECT 157.470 206.535 159.010 206.905 ;
        RECT 117.860 205.280 118.120 205.425 ;
        RECT 110.500 205.000 110.760 205.260 ;
        RECT 110.500 204.940 111.620 205.000 ;
        RECT 110.560 204.920 111.620 204.940 ;
        RECT 128.960 204.920 129.100 205.425 ;
        RECT 153.740 205.365 154.000 205.685 ;
        RECT 136.260 204.940 136.520 205.260 ;
        RECT 97.620 204.600 97.880 204.920 ;
        RECT 110.560 204.860 111.680 204.920 ;
        RECT 111.420 204.600 111.680 204.860 ;
        RECT 128.900 204.600 129.160 204.920 ;
        RECT 97.680 203.560 97.820 204.600 ;
        RECT 99.165 203.815 100.705 204.185 ;
        RECT 97.620 203.240 97.880 203.560 ;
        RECT 84.740 202.900 85.000 203.220 ;
        RECT 78.760 202.220 79.020 202.540 ;
        RECT 84.740 201.880 85.000 202.200 ;
        RECT 79.730 201.095 81.270 201.465 ;
        RECT 71.850 200.665 72.130 201.035 ;
        RECT 84.800 200.355 84.940 201.880 ;
        RECT 136.320 201.715 136.460 204.940 ;
        RECT 138.035 203.815 139.575 204.185 ;
        RECT 143.620 203.240 143.880 203.560 ;
        RECT 118.600 201.095 120.140 201.465 ;
        RECT 136.250 201.345 136.530 201.715 ;
        RECT 143.680 201.035 143.820 203.240 ;
        RECT 157.470 201.095 159.010 201.465 ;
        RECT 143.610 200.665 143.890 201.035 ;
        RECT 40.640 199.810 42.610 200.270 ;
        RECT 64.030 199.985 64.310 200.355 ;
        RECT 84.730 199.985 85.010 200.355 ;
        RECT 44.300 199.480 52.350 199.840 ;
        RECT 5.250 198.630 5.790 199.010 ;
        RECT 14.860 199.000 15.400 199.010 ;
        RECT 44.300 199.000 44.650 199.480 ;
        RECT 14.860 198.640 44.650 199.000 ;
        RECT 52.000 199.000 52.350 199.480 ;
        RECT 91.010 199.000 91.550 199.010 ;
        RECT 52.000 198.640 91.550 199.000 ;
        RECT 14.860 198.630 15.400 198.640 ;
        RECT 91.010 198.630 91.550 198.640 ;
        RECT 2.670 197.990 3.040 198.360 ;
        RECT 157.000 197.990 157.370 198.360 ;
        RECT 2.670 6.000 2.835 197.990 ;
        RECT 2.995 197.330 3.365 197.700 ;
        RECT 156.675 197.330 157.045 197.700 ;
        RECT 2.995 6.985 3.160 197.330 ;
        RECT 3.320 196.670 3.690 197.040 ;
        RECT 156.350 196.670 156.720 197.040 ;
        RECT 3.320 16.985 3.485 196.670 ;
        RECT 3.645 196.010 4.015 196.380 ;
        RECT 156.025 196.010 156.395 196.380 ;
        RECT 3.645 26.985 3.810 196.010 ;
        RECT 3.970 195.350 4.340 195.720 ;
        RECT 155.700 195.350 156.070 195.720 ;
        RECT 3.970 36.985 4.135 195.350 ;
        RECT 4.295 194.690 4.665 195.060 ;
        RECT 155.375 194.690 155.745 195.060 ;
        RECT 4.295 46.985 4.460 194.690 ;
        RECT 4.620 194.030 4.990 194.400 ;
        RECT 155.050 194.030 155.420 194.400 ;
        RECT 4.620 56.985 4.785 194.030 ;
        RECT 4.945 193.370 5.315 193.740 ;
        RECT 154.725 193.370 155.095 193.740 ;
        RECT 4.945 66.985 5.110 193.370 ;
        RECT 5.270 192.710 5.640 193.080 ;
        RECT 154.400 192.710 154.770 193.080 ;
        RECT 5.270 76.985 5.435 192.710 ;
        RECT 5.595 192.050 5.965 192.420 ;
        RECT 154.075 192.050 154.445 192.420 ;
        RECT 5.595 86.985 5.760 192.050 ;
        RECT 5.920 191.390 6.290 191.760 ;
        RECT 153.750 191.390 154.120 191.760 ;
        RECT 5.920 96.985 6.085 191.390 ;
        RECT 6.245 190.730 6.615 191.100 ;
        RECT 153.425 190.730 153.795 191.100 ;
        RECT 6.245 106.985 6.410 190.730 ;
        RECT 6.570 190.070 6.940 190.440 ;
        RECT 153.100 190.070 153.470 190.440 ;
        RECT 6.570 116.985 6.735 190.070 ;
        RECT 6.895 189.410 7.265 189.780 ;
        RECT 152.775 189.410 153.145 189.780 ;
        RECT 6.895 126.985 7.060 189.410 ;
        RECT 7.220 188.750 7.590 189.120 ;
        RECT 152.450 188.750 152.820 189.120 ;
        RECT 7.220 136.985 7.385 188.750 ;
        RECT 7.545 188.090 7.915 188.460 ;
        RECT 152.125 188.090 152.495 188.460 ;
        RECT 7.545 146.985 7.710 188.090 ;
        RECT 7.870 187.430 8.240 187.800 ;
        RECT 151.800 187.430 152.170 187.800 ;
        RECT 7.870 156.985 8.035 187.430 ;
        RECT 25.295 165.060 26.345 165.110 ;
        RECT 25.295 164.060 26.350 165.060 ;
        RECT 133.640 165.000 134.640 166.000 ;
        RECT 25.295 164.010 26.345 164.060 ;
        RECT 8.850 161.710 24.185 163.210 ;
        RECT 25.295 163.060 26.345 163.110 ;
        RECT 25.295 162.060 26.350 163.060 ;
        RECT 25.295 162.010 26.345 162.060 ;
        RECT 133.640 161.700 147.725 163.200 ;
        RECT 25.300 161.010 26.350 161.060 ;
        RECT 11.950 159.510 26.350 161.010 ;
        RECT 8.175 157.635 8.550 158.485 ;
        RECT 10.200 157.420 11.245 158.500 ;
        RECT 16.815 158.010 17.235 158.460 ;
        RECT 17.865 158.010 18.125 158.060 ;
        RECT 18.390 158.010 18.650 158.060 ;
        RECT 19.300 158.010 19.700 158.060 ;
        RECT 21.215 158.010 21.475 158.060 ;
        RECT 21.740 158.010 22.000 158.060 ;
        RECT 22.670 158.010 23.200 158.060 ;
        RECT 24.640 158.010 24.940 159.510 ;
        RECT 25.300 159.460 26.350 159.510 ;
        RECT 133.640 159.400 134.690 160.500 ;
        RECT 135.490 159.500 151.190 161.000 ;
        RECT 134.390 159.000 134.690 159.400 ;
        RECT 134.390 158.700 135.540 159.000 ;
        RECT 16.815 157.660 18.125 158.010 ;
        RECT 18.350 157.660 21.500 158.010 ;
        RECT 21.725 157.660 24.125 158.010 ;
        RECT 24.390 157.660 24.940 158.010 ;
        RECT 17.865 157.610 18.125 157.660 ;
        RECT 18.390 157.610 18.650 157.660 ;
        RECT 19.300 157.610 19.700 157.660 ;
        RECT 21.215 157.425 21.475 157.660 ;
        RECT 21.740 157.610 22.000 157.660 ;
        RECT 21.215 157.105 23.100 157.425 ;
        RECT 25.200 157.420 26.350 158.500 ;
        RECT 133.640 157.400 134.690 158.500 ;
        RECT 135.240 157.800 135.540 158.700 ;
        RECT 140.355 158.000 140.775 158.450 ;
        RECT 141.405 158.000 141.665 158.050 ;
        RECT 141.930 158.000 142.190 158.050 ;
        RECT 142.840 158.000 143.240 158.050 ;
        RECT 144.755 158.000 145.015 158.050 ;
        RECT 145.280 158.000 145.540 158.050 ;
        RECT 146.840 158.000 147.340 158.460 ;
        RECT 135.240 157.500 140.040 157.800 ;
        RECT 140.355 157.650 141.665 158.000 ;
        RECT 141.890 157.650 145.040 158.000 ;
        RECT 145.265 157.650 147.340 158.000 ;
        RECT 141.405 157.600 141.665 157.650 ;
        RECT 141.930 157.600 142.190 157.650 ;
        RECT 142.840 157.600 143.240 157.650 ;
        RECT 144.755 157.600 145.015 157.650 ;
        RECT 145.280 157.600 145.540 157.650 ;
        RECT 7.870 156.585 8.290 156.985 ;
        RECT 16.590 156.600 17.060 156.970 ;
        RECT 22.775 156.925 23.100 157.105 ;
        RECT 139.740 156.950 140.040 157.500 ;
        RECT 148.740 157.410 149.840 158.490 ;
        RECT 151.430 157.625 151.865 158.475 ;
        RECT 152.005 156.975 152.170 187.430 ;
        RECT 24.075 156.925 24.425 156.950 ;
        RECT 22.775 156.605 24.465 156.925 ;
        RECT 24.035 156.580 24.465 156.605 ;
        RECT 139.690 156.600 140.090 156.950 ;
        RECT 146.320 156.580 146.760 156.970 ;
        RECT 151.780 156.575 152.170 156.975 ;
        RECT 25.295 155.060 26.345 155.110 ;
        RECT 25.295 154.060 26.350 155.060 ;
        RECT 133.640 155.000 134.640 156.000 ;
        RECT 25.295 154.010 26.345 154.060 ;
        RECT 8.850 151.710 24.185 153.210 ;
        RECT 25.295 153.060 26.345 153.110 ;
        RECT 25.295 152.060 26.350 153.060 ;
        RECT 25.295 152.010 26.345 152.060 ;
        RECT 133.640 151.700 147.725 153.200 ;
        RECT 25.300 151.010 26.350 151.060 ;
        RECT 11.950 149.510 26.350 151.010 ;
        RECT 8.065 147.635 8.500 148.485 ;
        RECT 10.200 147.420 11.245 148.500 ;
        RECT 16.815 148.010 17.235 148.460 ;
        RECT 17.865 148.010 18.125 148.060 ;
        RECT 18.390 148.010 18.650 148.060 ;
        RECT 19.300 148.010 19.700 148.060 ;
        RECT 21.215 148.010 21.475 148.060 ;
        RECT 21.740 148.010 22.000 148.060 ;
        RECT 22.670 148.010 23.200 148.060 ;
        RECT 24.640 148.010 24.940 149.510 ;
        RECT 25.300 149.460 26.350 149.510 ;
        RECT 133.640 149.400 134.690 150.500 ;
        RECT 135.490 149.500 151.190 151.000 ;
        RECT 134.390 149.000 134.690 149.400 ;
        RECT 134.390 148.700 135.540 149.000 ;
        RECT 16.815 147.660 18.125 148.010 ;
        RECT 18.350 147.660 21.500 148.010 ;
        RECT 21.725 147.660 24.125 148.010 ;
        RECT 24.390 147.660 24.940 148.010 ;
        RECT 17.865 147.610 18.125 147.660 ;
        RECT 18.390 147.610 18.650 147.660 ;
        RECT 19.300 147.610 19.700 147.660 ;
        RECT 21.215 147.425 21.475 147.660 ;
        RECT 21.740 147.610 22.000 147.660 ;
        RECT 21.215 147.105 23.100 147.425 ;
        RECT 25.200 147.420 26.350 148.500 ;
        RECT 133.640 147.400 134.690 148.500 ;
        RECT 135.240 147.800 135.540 148.700 ;
        RECT 140.355 148.000 140.775 148.450 ;
        RECT 141.405 148.000 141.665 148.050 ;
        RECT 141.930 148.000 142.190 148.050 ;
        RECT 142.840 148.000 143.240 148.050 ;
        RECT 144.755 148.000 145.015 148.050 ;
        RECT 145.280 148.000 145.540 148.050 ;
        RECT 146.840 148.000 147.340 148.460 ;
        RECT 135.240 147.500 140.040 147.800 ;
        RECT 140.355 147.650 141.665 148.000 ;
        RECT 141.890 147.650 145.040 148.000 ;
        RECT 145.265 147.650 147.340 148.000 ;
        RECT 141.405 147.600 141.665 147.650 ;
        RECT 141.930 147.600 142.190 147.650 ;
        RECT 142.840 147.600 143.240 147.650 ;
        RECT 144.755 147.600 145.015 147.650 ;
        RECT 145.280 147.600 145.540 147.650 ;
        RECT 7.545 146.585 7.925 146.985 ;
        RECT 16.590 146.600 17.060 146.970 ;
        RECT 22.775 146.925 23.100 147.105 ;
        RECT 139.740 146.950 140.040 147.500 ;
        RECT 148.740 147.410 149.840 148.490 ;
        RECT 151.540 147.625 151.975 148.475 ;
        RECT 152.330 146.975 152.495 188.090 ;
        RECT 24.075 146.925 24.425 146.950 ;
        RECT 22.775 146.605 24.465 146.925 ;
        RECT 24.035 146.580 24.465 146.605 ;
        RECT 139.690 146.600 140.090 146.950 ;
        RECT 146.320 146.580 146.760 146.970 ;
        RECT 152.115 146.575 152.495 146.975 ;
        RECT 25.295 145.060 26.345 145.110 ;
        RECT 25.295 144.060 26.350 145.060 ;
        RECT 133.640 145.000 134.640 146.000 ;
        RECT 25.295 144.010 26.345 144.060 ;
        RECT 8.850 141.710 24.185 143.210 ;
        RECT 25.295 143.060 26.345 143.110 ;
        RECT 25.295 142.060 26.350 143.060 ;
        RECT 25.295 142.010 26.345 142.060 ;
        RECT 133.640 141.700 147.725 143.200 ;
        RECT 25.300 141.010 26.350 141.060 ;
        RECT 11.950 139.510 26.350 141.010 ;
        RECT 8.065 137.635 8.500 138.485 ;
        RECT 10.200 137.420 11.245 138.500 ;
        RECT 16.815 138.010 17.235 138.460 ;
        RECT 17.865 138.010 18.125 138.060 ;
        RECT 18.390 138.010 18.650 138.060 ;
        RECT 19.300 138.010 19.700 138.060 ;
        RECT 21.215 138.010 21.475 138.060 ;
        RECT 21.740 138.010 22.000 138.060 ;
        RECT 22.670 138.010 23.200 138.060 ;
        RECT 24.640 138.010 24.940 139.510 ;
        RECT 25.300 139.460 26.350 139.510 ;
        RECT 133.640 139.400 134.690 140.500 ;
        RECT 135.490 139.500 151.190 141.000 ;
        RECT 134.390 139.000 134.690 139.400 ;
        RECT 134.390 138.700 135.540 139.000 ;
        RECT 16.815 137.660 18.125 138.010 ;
        RECT 18.350 137.660 21.500 138.010 ;
        RECT 21.725 137.660 24.125 138.010 ;
        RECT 24.390 137.660 24.940 138.010 ;
        RECT 17.865 137.610 18.125 137.660 ;
        RECT 18.390 137.610 18.650 137.660 ;
        RECT 19.300 137.610 19.700 137.660 ;
        RECT 21.215 137.425 21.475 137.660 ;
        RECT 21.740 137.610 22.000 137.660 ;
        RECT 21.215 137.105 23.100 137.425 ;
        RECT 25.200 137.420 26.350 138.500 ;
        RECT 133.640 137.400 134.690 138.500 ;
        RECT 135.240 137.800 135.540 138.700 ;
        RECT 140.355 138.000 140.775 138.450 ;
        RECT 141.405 138.000 141.665 138.050 ;
        RECT 141.930 138.000 142.190 138.050 ;
        RECT 142.840 138.000 143.240 138.050 ;
        RECT 144.755 138.000 145.015 138.050 ;
        RECT 145.280 138.000 145.540 138.050 ;
        RECT 146.840 138.000 147.340 138.460 ;
        RECT 135.240 137.500 140.040 137.800 ;
        RECT 140.355 137.650 141.665 138.000 ;
        RECT 141.890 137.650 145.040 138.000 ;
        RECT 145.265 137.650 147.340 138.000 ;
        RECT 141.405 137.600 141.665 137.650 ;
        RECT 141.930 137.600 142.190 137.650 ;
        RECT 142.840 137.600 143.240 137.650 ;
        RECT 144.755 137.600 145.015 137.650 ;
        RECT 145.280 137.600 145.540 137.650 ;
        RECT 7.220 136.585 7.645 136.985 ;
        RECT 16.590 136.600 17.060 136.970 ;
        RECT 22.775 136.925 23.100 137.105 ;
        RECT 139.740 136.950 140.040 137.500 ;
        RECT 148.740 137.410 149.840 138.490 ;
        RECT 151.540 137.625 151.975 138.475 ;
        RECT 152.655 136.975 152.820 188.750 ;
        RECT 24.075 136.925 24.425 136.950 ;
        RECT 22.775 136.605 24.465 136.925 ;
        RECT 24.035 136.580 24.465 136.605 ;
        RECT 139.690 136.600 140.090 136.950 ;
        RECT 146.320 136.580 146.760 136.970 ;
        RECT 152.440 136.575 152.820 136.975 ;
        RECT 25.295 135.060 26.345 135.110 ;
        RECT 25.295 134.060 26.350 135.060 ;
        RECT 133.640 135.000 134.640 136.000 ;
        RECT 25.295 134.010 26.345 134.060 ;
        RECT 8.850 131.710 24.185 133.210 ;
        RECT 25.295 133.060 26.345 133.110 ;
        RECT 25.295 132.060 26.350 133.060 ;
        RECT 25.295 132.010 26.345 132.060 ;
        RECT 133.640 131.700 147.725 133.200 ;
        RECT 25.300 131.010 26.350 131.060 ;
        RECT 11.950 129.510 26.350 131.010 ;
        RECT 8.065 127.635 8.500 128.485 ;
        RECT 10.200 127.420 11.245 128.500 ;
        RECT 16.815 128.010 17.235 128.460 ;
        RECT 17.865 128.010 18.125 128.060 ;
        RECT 18.390 128.010 18.650 128.060 ;
        RECT 19.300 128.010 19.700 128.060 ;
        RECT 21.215 128.010 21.475 128.060 ;
        RECT 21.740 128.010 22.000 128.060 ;
        RECT 22.670 128.010 23.200 128.060 ;
        RECT 24.640 128.010 24.940 129.510 ;
        RECT 25.300 129.460 26.350 129.510 ;
        RECT 133.640 129.400 134.690 130.500 ;
        RECT 135.490 129.500 151.190 131.000 ;
        RECT 134.390 129.000 134.690 129.400 ;
        RECT 134.390 128.700 135.540 129.000 ;
        RECT 16.815 127.660 18.125 128.010 ;
        RECT 18.350 127.660 21.500 128.010 ;
        RECT 21.725 127.660 24.125 128.010 ;
        RECT 24.390 127.660 24.940 128.010 ;
        RECT 17.865 127.610 18.125 127.660 ;
        RECT 18.390 127.610 18.650 127.660 ;
        RECT 19.300 127.610 19.700 127.660 ;
        RECT 21.215 127.425 21.475 127.660 ;
        RECT 21.740 127.610 22.000 127.660 ;
        RECT 21.215 127.105 23.100 127.425 ;
        RECT 25.200 127.420 26.350 128.500 ;
        RECT 133.640 127.400 134.690 128.500 ;
        RECT 135.240 127.800 135.540 128.700 ;
        RECT 140.355 128.000 140.775 128.450 ;
        RECT 141.405 128.000 141.665 128.050 ;
        RECT 141.930 128.000 142.190 128.050 ;
        RECT 142.840 128.000 143.240 128.050 ;
        RECT 144.755 128.000 145.015 128.050 ;
        RECT 145.280 128.000 145.540 128.050 ;
        RECT 146.840 128.000 147.340 128.460 ;
        RECT 135.240 127.500 140.040 127.800 ;
        RECT 140.355 127.650 141.665 128.000 ;
        RECT 141.890 127.650 145.040 128.000 ;
        RECT 145.265 127.650 147.340 128.000 ;
        RECT 141.405 127.600 141.665 127.650 ;
        RECT 141.930 127.600 142.190 127.650 ;
        RECT 142.840 127.600 143.240 127.650 ;
        RECT 144.755 127.600 145.015 127.650 ;
        RECT 145.280 127.600 145.540 127.650 ;
        RECT 6.895 126.585 7.320 126.985 ;
        RECT 16.590 126.600 17.060 126.970 ;
        RECT 22.775 126.925 23.100 127.105 ;
        RECT 139.740 126.950 140.040 127.500 ;
        RECT 148.740 127.410 149.840 128.490 ;
        RECT 151.540 127.625 151.975 128.475 ;
        RECT 152.980 126.975 153.145 189.410 ;
        RECT 24.075 126.925 24.425 126.950 ;
        RECT 22.775 126.605 24.465 126.925 ;
        RECT 24.035 126.580 24.465 126.605 ;
        RECT 139.690 126.600 140.090 126.950 ;
        RECT 146.320 126.580 146.760 126.970 ;
        RECT 152.765 126.575 153.145 126.975 ;
        RECT 25.295 125.060 26.345 125.110 ;
        RECT 25.295 124.060 26.350 125.060 ;
        RECT 133.640 125.000 134.640 126.000 ;
        RECT 25.295 124.010 26.345 124.060 ;
        RECT 8.850 121.710 24.185 123.210 ;
        RECT 25.295 123.060 26.345 123.110 ;
        RECT 25.295 122.060 26.350 123.060 ;
        RECT 25.295 122.010 26.345 122.060 ;
        RECT 133.640 121.700 147.725 123.200 ;
        RECT 25.300 121.010 26.350 121.060 ;
        RECT 11.950 119.510 26.350 121.010 ;
        RECT 8.065 117.635 8.500 118.485 ;
        RECT 10.200 117.420 11.245 118.500 ;
        RECT 16.815 118.010 17.235 118.460 ;
        RECT 17.865 118.010 18.125 118.060 ;
        RECT 18.390 118.010 18.650 118.060 ;
        RECT 19.300 118.010 19.700 118.060 ;
        RECT 21.215 118.010 21.475 118.060 ;
        RECT 21.740 118.010 22.000 118.060 ;
        RECT 22.670 118.010 23.200 118.060 ;
        RECT 24.640 118.010 24.940 119.510 ;
        RECT 25.300 119.460 26.350 119.510 ;
        RECT 133.640 119.400 134.690 120.500 ;
        RECT 135.490 119.500 151.190 121.000 ;
        RECT 134.390 119.000 134.690 119.400 ;
        RECT 134.390 118.700 135.540 119.000 ;
        RECT 16.815 117.660 18.125 118.010 ;
        RECT 18.350 117.660 21.500 118.010 ;
        RECT 21.725 117.660 24.125 118.010 ;
        RECT 24.390 117.660 24.940 118.010 ;
        RECT 17.865 117.610 18.125 117.660 ;
        RECT 18.390 117.610 18.650 117.660 ;
        RECT 19.300 117.610 19.700 117.660 ;
        RECT 21.215 117.425 21.475 117.660 ;
        RECT 21.740 117.610 22.000 117.660 ;
        RECT 21.215 117.105 23.100 117.425 ;
        RECT 25.200 117.420 26.350 118.500 ;
        RECT 133.640 117.400 134.690 118.500 ;
        RECT 135.240 117.800 135.540 118.700 ;
        RECT 140.355 118.000 140.775 118.450 ;
        RECT 141.405 118.000 141.665 118.050 ;
        RECT 141.930 118.000 142.190 118.050 ;
        RECT 142.840 118.000 143.240 118.050 ;
        RECT 144.755 118.000 145.015 118.050 ;
        RECT 145.280 118.000 145.540 118.050 ;
        RECT 146.840 118.000 147.340 118.460 ;
        RECT 135.240 117.500 140.040 117.800 ;
        RECT 140.355 117.650 141.665 118.000 ;
        RECT 141.890 117.650 145.040 118.000 ;
        RECT 145.265 117.650 147.340 118.000 ;
        RECT 141.405 117.600 141.665 117.650 ;
        RECT 141.930 117.600 142.190 117.650 ;
        RECT 142.840 117.600 143.240 117.650 ;
        RECT 144.755 117.600 145.015 117.650 ;
        RECT 145.280 117.600 145.540 117.650 ;
        RECT 6.570 116.585 6.950 116.985 ;
        RECT 16.590 116.600 17.060 116.970 ;
        RECT 22.775 116.925 23.100 117.105 ;
        RECT 139.740 116.950 140.040 117.500 ;
        RECT 148.740 117.410 149.840 118.490 ;
        RECT 151.540 117.625 151.975 118.475 ;
        RECT 153.305 116.975 153.470 190.070 ;
        RECT 24.075 116.925 24.425 116.950 ;
        RECT 22.775 116.605 24.465 116.925 ;
        RECT 24.035 116.580 24.465 116.605 ;
        RECT 139.690 116.600 140.090 116.950 ;
        RECT 146.320 116.580 146.760 116.970 ;
        RECT 153.090 116.575 153.470 116.975 ;
        RECT 25.295 115.060 26.345 115.110 ;
        RECT 25.295 114.060 26.350 115.060 ;
        RECT 133.640 115.000 134.640 116.000 ;
        RECT 25.295 114.010 26.345 114.060 ;
        RECT 8.850 111.710 24.185 113.210 ;
        RECT 25.295 113.060 26.345 113.110 ;
        RECT 25.295 112.060 26.350 113.060 ;
        RECT 25.295 112.010 26.345 112.060 ;
        RECT 133.640 111.700 147.725 113.200 ;
        RECT 25.300 111.010 26.350 111.060 ;
        RECT 11.950 109.510 26.350 111.010 ;
        RECT 8.065 107.635 8.500 108.485 ;
        RECT 10.200 107.420 11.245 108.500 ;
        RECT 16.815 108.010 17.235 108.460 ;
        RECT 17.865 108.010 18.125 108.060 ;
        RECT 18.390 108.010 18.650 108.060 ;
        RECT 19.300 108.010 19.700 108.060 ;
        RECT 21.215 108.010 21.475 108.060 ;
        RECT 21.740 108.010 22.000 108.060 ;
        RECT 22.670 108.010 23.200 108.060 ;
        RECT 24.640 108.010 24.940 109.510 ;
        RECT 25.300 109.460 26.350 109.510 ;
        RECT 133.640 109.400 134.690 110.500 ;
        RECT 135.490 109.500 151.190 111.000 ;
        RECT 134.390 109.000 134.690 109.400 ;
        RECT 134.390 108.700 135.540 109.000 ;
        RECT 16.815 107.660 18.125 108.010 ;
        RECT 18.350 107.660 21.500 108.010 ;
        RECT 21.725 107.660 24.125 108.010 ;
        RECT 24.390 107.660 24.940 108.010 ;
        RECT 17.865 107.610 18.125 107.660 ;
        RECT 18.390 107.610 18.650 107.660 ;
        RECT 19.300 107.610 19.700 107.660 ;
        RECT 21.215 107.425 21.475 107.660 ;
        RECT 21.740 107.610 22.000 107.660 ;
        RECT 21.215 107.105 23.100 107.425 ;
        RECT 25.200 107.420 26.350 108.500 ;
        RECT 133.640 107.400 134.690 108.500 ;
        RECT 135.240 107.800 135.540 108.700 ;
        RECT 140.355 108.000 140.775 108.450 ;
        RECT 141.405 108.000 141.665 108.050 ;
        RECT 141.930 108.000 142.190 108.050 ;
        RECT 142.840 108.000 143.240 108.050 ;
        RECT 144.755 108.000 145.015 108.050 ;
        RECT 145.280 108.000 145.540 108.050 ;
        RECT 146.840 108.000 147.340 108.460 ;
        RECT 135.240 107.500 140.040 107.800 ;
        RECT 140.355 107.650 141.665 108.000 ;
        RECT 141.890 107.650 145.040 108.000 ;
        RECT 145.265 107.650 147.340 108.000 ;
        RECT 141.405 107.600 141.665 107.650 ;
        RECT 141.930 107.600 142.190 107.650 ;
        RECT 142.840 107.600 143.240 107.650 ;
        RECT 144.755 107.600 145.015 107.650 ;
        RECT 145.280 107.600 145.540 107.650 ;
        RECT 6.245 106.585 6.670 106.985 ;
        RECT 16.590 106.600 17.060 106.970 ;
        RECT 22.775 106.925 23.100 107.105 ;
        RECT 139.740 106.950 140.040 107.500 ;
        RECT 148.740 107.410 149.840 108.490 ;
        RECT 151.540 107.625 151.975 108.475 ;
        RECT 153.630 106.975 153.795 190.730 ;
        RECT 24.075 106.925 24.425 106.950 ;
        RECT 22.775 106.605 24.465 106.925 ;
        RECT 24.035 106.580 24.465 106.605 ;
        RECT 139.690 106.600 140.090 106.950 ;
        RECT 146.320 106.580 146.760 106.970 ;
        RECT 153.415 106.575 153.795 106.975 ;
        RECT 25.295 105.060 26.345 105.110 ;
        RECT 25.295 104.060 26.350 105.060 ;
        RECT 133.640 105.000 134.640 106.000 ;
        RECT 25.295 104.010 26.345 104.060 ;
        RECT 8.850 101.710 24.185 103.210 ;
        RECT 25.295 103.060 26.345 103.110 ;
        RECT 25.295 102.060 26.350 103.060 ;
        RECT 25.295 102.010 26.345 102.060 ;
        RECT 133.640 101.700 147.725 103.200 ;
        RECT 25.300 101.010 26.350 101.060 ;
        RECT 11.950 99.510 26.350 101.010 ;
        RECT 8.065 97.635 8.500 98.485 ;
        RECT 10.200 97.420 11.245 98.500 ;
        RECT 16.815 98.010 17.235 98.460 ;
        RECT 17.865 98.010 18.125 98.060 ;
        RECT 18.390 98.010 18.650 98.060 ;
        RECT 19.300 98.010 19.700 98.060 ;
        RECT 21.215 98.010 21.475 98.060 ;
        RECT 21.740 98.010 22.000 98.060 ;
        RECT 22.670 98.010 23.200 98.060 ;
        RECT 24.640 98.010 24.940 99.510 ;
        RECT 25.300 99.460 26.350 99.510 ;
        RECT 133.640 99.400 134.690 100.500 ;
        RECT 135.490 99.500 151.190 101.000 ;
        RECT 134.390 99.000 134.690 99.400 ;
        RECT 134.390 98.700 135.540 99.000 ;
        RECT 16.815 97.660 18.125 98.010 ;
        RECT 18.350 97.660 21.500 98.010 ;
        RECT 21.725 97.660 24.125 98.010 ;
        RECT 24.390 97.660 24.940 98.010 ;
        RECT 17.865 97.610 18.125 97.660 ;
        RECT 18.390 97.610 18.650 97.660 ;
        RECT 19.300 97.610 19.700 97.660 ;
        RECT 21.215 97.425 21.475 97.660 ;
        RECT 21.740 97.610 22.000 97.660 ;
        RECT 21.215 97.105 23.100 97.425 ;
        RECT 25.200 97.420 26.350 98.500 ;
        RECT 133.640 97.400 134.690 98.500 ;
        RECT 135.240 97.800 135.540 98.700 ;
        RECT 140.355 98.000 140.775 98.450 ;
        RECT 141.405 98.000 141.665 98.050 ;
        RECT 141.930 98.000 142.190 98.050 ;
        RECT 142.840 98.000 143.240 98.050 ;
        RECT 144.755 98.000 145.015 98.050 ;
        RECT 145.280 98.000 145.540 98.050 ;
        RECT 146.840 98.000 147.340 98.460 ;
        RECT 135.240 97.500 140.040 97.800 ;
        RECT 140.355 97.650 141.665 98.000 ;
        RECT 141.890 97.650 145.040 98.000 ;
        RECT 145.265 97.650 147.340 98.000 ;
        RECT 141.405 97.600 141.665 97.650 ;
        RECT 141.930 97.600 142.190 97.650 ;
        RECT 142.840 97.600 143.240 97.650 ;
        RECT 144.755 97.600 145.015 97.650 ;
        RECT 145.280 97.600 145.540 97.650 ;
        RECT 5.920 96.585 6.300 96.985 ;
        RECT 16.590 96.600 17.060 96.970 ;
        RECT 22.775 96.925 23.100 97.105 ;
        RECT 139.740 96.950 140.040 97.500 ;
        RECT 148.740 97.410 149.840 98.490 ;
        RECT 151.540 97.625 151.975 98.475 ;
        RECT 153.955 96.975 154.120 191.390 ;
        RECT 24.075 96.925 24.425 96.950 ;
        RECT 22.775 96.605 24.465 96.925 ;
        RECT 24.035 96.580 24.465 96.605 ;
        RECT 139.690 96.600 140.090 96.950 ;
        RECT 146.320 96.580 146.760 96.970 ;
        RECT 153.740 96.575 154.120 96.975 ;
        RECT 25.295 95.060 26.345 95.110 ;
        RECT 25.295 94.060 26.350 95.060 ;
        RECT 133.640 95.000 134.640 96.000 ;
        RECT 25.295 94.010 26.345 94.060 ;
        RECT 8.850 91.710 24.185 93.210 ;
        RECT 25.295 93.060 26.345 93.110 ;
        RECT 25.295 92.060 26.350 93.060 ;
        RECT 25.295 92.010 26.345 92.060 ;
        RECT 133.640 91.700 147.725 93.200 ;
        RECT 25.300 91.010 26.350 91.060 ;
        RECT 11.950 89.510 26.350 91.010 ;
        RECT 8.065 87.635 8.500 88.485 ;
        RECT 10.200 87.420 11.245 88.500 ;
        RECT 16.815 88.010 17.235 88.460 ;
        RECT 17.865 88.010 18.125 88.060 ;
        RECT 18.390 88.010 18.650 88.060 ;
        RECT 19.300 88.010 19.700 88.060 ;
        RECT 21.215 88.010 21.475 88.060 ;
        RECT 21.740 88.010 22.000 88.060 ;
        RECT 22.670 88.010 23.200 88.060 ;
        RECT 24.640 88.010 24.940 89.510 ;
        RECT 25.300 89.460 26.350 89.510 ;
        RECT 133.640 89.400 134.690 90.500 ;
        RECT 135.490 89.500 151.190 91.000 ;
        RECT 134.390 89.000 134.690 89.400 ;
        RECT 134.390 88.700 135.540 89.000 ;
        RECT 16.815 87.660 18.125 88.010 ;
        RECT 18.350 87.660 21.500 88.010 ;
        RECT 21.725 87.660 24.125 88.010 ;
        RECT 24.390 87.660 24.940 88.010 ;
        RECT 17.865 87.610 18.125 87.660 ;
        RECT 18.390 87.610 18.650 87.660 ;
        RECT 19.300 87.610 19.700 87.660 ;
        RECT 21.215 87.425 21.475 87.660 ;
        RECT 21.740 87.610 22.000 87.660 ;
        RECT 21.215 87.105 23.100 87.425 ;
        RECT 25.200 87.420 26.350 88.500 ;
        RECT 133.640 87.400 134.690 88.500 ;
        RECT 135.240 87.800 135.540 88.700 ;
        RECT 140.355 88.000 140.775 88.450 ;
        RECT 141.405 88.000 141.665 88.050 ;
        RECT 141.930 88.000 142.190 88.050 ;
        RECT 142.840 88.000 143.240 88.050 ;
        RECT 144.755 88.000 145.015 88.050 ;
        RECT 145.280 88.000 145.540 88.050 ;
        RECT 146.840 88.000 147.340 88.460 ;
        RECT 135.240 87.500 140.040 87.800 ;
        RECT 140.355 87.650 141.665 88.000 ;
        RECT 141.890 87.650 145.040 88.000 ;
        RECT 145.265 87.650 147.340 88.000 ;
        RECT 141.405 87.600 141.665 87.650 ;
        RECT 141.930 87.600 142.190 87.650 ;
        RECT 142.840 87.600 143.240 87.650 ;
        RECT 144.755 87.600 145.015 87.650 ;
        RECT 145.280 87.600 145.540 87.650 ;
        RECT 5.595 86.585 5.975 86.985 ;
        RECT 16.590 86.600 17.060 86.970 ;
        RECT 22.775 86.925 23.100 87.105 ;
        RECT 139.740 86.950 140.040 87.500 ;
        RECT 148.740 87.410 149.840 88.490 ;
        RECT 151.540 87.625 151.975 88.475 ;
        RECT 154.280 86.975 154.445 192.050 ;
        RECT 24.075 86.925 24.425 86.950 ;
        RECT 22.775 86.605 24.465 86.925 ;
        RECT 24.035 86.580 24.465 86.605 ;
        RECT 139.690 86.600 140.090 86.950 ;
        RECT 146.320 86.580 146.760 86.970 ;
        RECT 154.065 86.575 154.445 86.975 ;
        RECT 25.295 85.060 26.345 85.110 ;
        RECT 25.295 84.060 26.350 85.060 ;
        RECT 133.640 85.000 134.640 86.000 ;
        RECT 25.295 84.010 26.345 84.060 ;
        RECT 8.850 81.710 24.185 83.210 ;
        RECT 25.295 83.060 26.345 83.110 ;
        RECT 25.295 82.060 26.350 83.060 ;
        RECT 25.295 82.010 26.345 82.060 ;
        RECT 133.640 81.700 147.725 83.200 ;
        RECT 25.300 81.010 26.350 81.060 ;
        RECT 11.950 79.510 26.350 81.010 ;
        RECT 8.065 77.635 8.500 78.485 ;
        RECT 10.200 77.420 11.245 78.500 ;
        RECT 16.815 78.010 17.235 78.460 ;
        RECT 17.865 78.010 18.125 78.060 ;
        RECT 18.390 78.010 18.650 78.060 ;
        RECT 19.300 78.010 19.700 78.060 ;
        RECT 21.215 78.010 21.475 78.060 ;
        RECT 21.740 78.010 22.000 78.060 ;
        RECT 22.670 78.010 23.200 78.060 ;
        RECT 24.640 78.010 24.940 79.510 ;
        RECT 25.300 79.460 26.350 79.510 ;
        RECT 133.640 79.400 134.690 80.500 ;
        RECT 135.490 79.500 151.190 81.000 ;
        RECT 134.390 79.000 134.690 79.400 ;
        RECT 134.390 78.700 135.540 79.000 ;
        RECT 16.815 77.660 18.125 78.010 ;
        RECT 18.350 77.660 21.500 78.010 ;
        RECT 21.725 77.660 24.125 78.010 ;
        RECT 24.390 77.660 24.940 78.010 ;
        RECT 17.865 77.610 18.125 77.660 ;
        RECT 18.390 77.610 18.650 77.660 ;
        RECT 19.300 77.610 19.700 77.660 ;
        RECT 21.215 77.425 21.475 77.660 ;
        RECT 21.740 77.610 22.000 77.660 ;
        RECT 21.215 77.105 23.100 77.425 ;
        RECT 25.200 77.420 26.350 78.500 ;
        RECT 133.640 77.400 134.690 78.500 ;
        RECT 135.240 77.800 135.540 78.700 ;
        RECT 140.355 78.000 140.775 78.450 ;
        RECT 141.405 78.000 141.665 78.050 ;
        RECT 141.930 78.000 142.190 78.050 ;
        RECT 142.840 78.000 143.240 78.050 ;
        RECT 144.755 78.000 145.015 78.050 ;
        RECT 145.280 78.000 145.540 78.050 ;
        RECT 146.840 78.000 147.340 78.460 ;
        RECT 135.240 77.500 140.040 77.800 ;
        RECT 140.355 77.650 141.665 78.000 ;
        RECT 141.890 77.650 145.040 78.000 ;
        RECT 145.265 77.650 147.340 78.000 ;
        RECT 141.405 77.600 141.665 77.650 ;
        RECT 141.930 77.600 142.190 77.650 ;
        RECT 142.840 77.600 143.240 77.650 ;
        RECT 144.755 77.600 145.015 77.650 ;
        RECT 145.280 77.600 145.540 77.650 ;
        RECT 5.270 76.585 5.650 76.985 ;
        RECT 16.590 76.600 17.060 76.970 ;
        RECT 22.775 76.925 23.100 77.105 ;
        RECT 139.740 76.950 140.040 77.500 ;
        RECT 148.740 77.410 149.840 78.490 ;
        RECT 151.540 77.625 151.975 78.475 ;
        RECT 154.605 76.975 154.770 192.710 ;
        RECT 24.075 76.925 24.425 76.950 ;
        RECT 22.775 76.605 24.465 76.925 ;
        RECT 24.035 76.580 24.465 76.605 ;
        RECT 139.690 76.600 140.090 76.950 ;
        RECT 146.320 76.580 146.760 76.970 ;
        RECT 154.390 76.575 154.770 76.975 ;
        RECT 25.295 75.060 26.345 75.110 ;
        RECT 25.295 74.060 26.350 75.060 ;
        RECT 133.640 75.000 134.640 76.000 ;
        RECT 25.295 74.010 26.345 74.060 ;
        RECT 8.850 71.710 24.185 73.210 ;
        RECT 25.295 73.060 26.345 73.110 ;
        RECT 25.295 72.060 26.350 73.060 ;
        RECT 25.295 72.010 26.345 72.060 ;
        RECT 133.640 71.700 147.725 73.200 ;
        RECT 25.300 71.010 26.350 71.060 ;
        RECT 11.950 69.510 26.350 71.010 ;
        RECT 8.065 67.635 8.500 68.485 ;
        RECT 10.200 67.420 11.245 68.500 ;
        RECT 16.815 68.010 17.235 68.460 ;
        RECT 17.865 68.010 18.125 68.060 ;
        RECT 18.390 68.010 18.650 68.060 ;
        RECT 19.300 68.010 19.700 68.060 ;
        RECT 21.215 68.010 21.475 68.060 ;
        RECT 21.740 68.010 22.000 68.060 ;
        RECT 22.670 68.010 23.200 68.060 ;
        RECT 24.640 68.010 24.940 69.510 ;
        RECT 25.300 69.460 26.350 69.510 ;
        RECT 133.640 69.400 134.690 70.500 ;
        RECT 135.490 69.500 151.190 71.000 ;
        RECT 134.390 69.000 134.690 69.400 ;
        RECT 134.390 68.700 135.540 69.000 ;
        RECT 16.815 67.660 18.125 68.010 ;
        RECT 18.350 67.660 21.500 68.010 ;
        RECT 21.725 67.660 24.125 68.010 ;
        RECT 24.390 67.660 24.940 68.010 ;
        RECT 17.865 67.610 18.125 67.660 ;
        RECT 18.390 67.610 18.650 67.660 ;
        RECT 19.300 67.610 19.700 67.660 ;
        RECT 21.215 67.425 21.475 67.660 ;
        RECT 21.740 67.610 22.000 67.660 ;
        RECT 21.215 67.105 23.100 67.425 ;
        RECT 25.200 67.420 26.350 68.500 ;
        RECT 133.640 67.400 134.690 68.500 ;
        RECT 135.240 67.800 135.540 68.700 ;
        RECT 140.355 68.000 140.775 68.450 ;
        RECT 141.405 68.000 141.665 68.050 ;
        RECT 141.930 68.000 142.190 68.050 ;
        RECT 142.840 68.000 143.240 68.050 ;
        RECT 144.755 68.000 145.015 68.050 ;
        RECT 145.280 68.000 145.540 68.050 ;
        RECT 146.840 68.000 147.340 68.460 ;
        RECT 135.240 67.500 140.040 67.800 ;
        RECT 140.355 67.650 141.665 68.000 ;
        RECT 141.890 67.650 145.040 68.000 ;
        RECT 145.265 67.650 147.340 68.000 ;
        RECT 141.405 67.600 141.665 67.650 ;
        RECT 141.930 67.600 142.190 67.650 ;
        RECT 142.840 67.600 143.240 67.650 ;
        RECT 144.755 67.600 145.015 67.650 ;
        RECT 145.280 67.600 145.540 67.650 ;
        RECT 4.945 66.585 5.325 66.985 ;
        RECT 16.590 66.600 17.060 66.970 ;
        RECT 22.775 66.925 23.100 67.105 ;
        RECT 139.740 66.950 140.040 67.500 ;
        RECT 148.740 67.410 149.840 68.490 ;
        RECT 151.540 67.625 151.975 68.475 ;
        RECT 154.930 66.975 155.095 193.370 ;
        RECT 24.075 66.925 24.425 66.950 ;
        RECT 22.775 66.605 24.465 66.925 ;
        RECT 24.035 66.580 24.465 66.605 ;
        RECT 139.690 66.600 140.090 66.950 ;
        RECT 146.320 66.580 146.760 66.970 ;
        RECT 154.715 66.575 155.095 66.975 ;
        RECT 25.295 65.060 26.345 65.110 ;
        RECT 25.295 64.060 26.350 65.060 ;
        RECT 133.640 65.000 134.640 66.000 ;
        RECT 25.295 64.010 26.345 64.060 ;
        RECT 8.850 61.710 24.185 63.210 ;
        RECT 25.295 63.060 26.345 63.110 ;
        RECT 25.295 62.060 26.350 63.060 ;
        RECT 25.295 62.010 26.345 62.060 ;
        RECT 133.640 61.700 147.725 63.200 ;
        RECT 25.300 61.010 26.350 61.060 ;
        RECT 11.950 59.510 26.350 61.010 ;
        RECT 8.065 57.635 8.500 58.485 ;
        RECT 10.200 57.420 11.245 58.500 ;
        RECT 16.815 58.010 17.235 58.460 ;
        RECT 17.865 58.010 18.125 58.060 ;
        RECT 18.390 58.010 18.650 58.060 ;
        RECT 19.300 58.010 19.700 58.060 ;
        RECT 21.215 58.010 21.475 58.060 ;
        RECT 21.740 58.010 22.000 58.060 ;
        RECT 22.670 58.010 23.200 58.060 ;
        RECT 24.640 58.010 24.940 59.510 ;
        RECT 25.300 59.460 26.350 59.510 ;
        RECT 133.640 59.400 134.690 60.500 ;
        RECT 135.490 59.500 151.190 61.000 ;
        RECT 134.390 59.000 134.690 59.400 ;
        RECT 134.390 58.700 135.540 59.000 ;
        RECT 16.815 57.660 18.125 58.010 ;
        RECT 18.350 57.660 21.500 58.010 ;
        RECT 21.725 57.660 24.125 58.010 ;
        RECT 24.390 57.660 24.940 58.010 ;
        RECT 17.865 57.610 18.125 57.660 ;
        RECT 18.390 57.610 18.650 57.660 ;
        RECT 19.300 57.610 19.700 57.660 ;
        RECT 21.215 57.425 21.475 57.660 ;
        RECT 21.740 57.610 22.000 57.660 ;
        RECT 21.215 57.105 23.100 57.425 ;
        RECT 25.200 57.420 26.350 58.500 ;
        RECT 133.640 57.400 134.690 58.500 ;
        RECT 135.240 57.800 135.540 58.700 ;
        RECT 140.355 58.000 140.775 58.450 ;
        RECT 141.405 58.000 141.665 58.050 ;
        RECT 141.930 58.000 142.190 58.050 ;
        RECT 142.840 58.000 143.240 58.050 ;
        RECT 144.755 58.000 145.015 58.050 ;
        RECT 145.280 58.000 145.540 58.050 ;
        RECT 146.840 58.000 147.340 58.460 ;
        RECT 135.240 57.500 140.040 57.800 ;
        RECT 140.355 57.650 141.665 58.000 ;
        RECT 141.890 57.650 145.040 58.000 ;
        RECT 145.265 57.650 147.340 58.000 ;
        RECT 141.405 57.600 141.665 57.650 ;
        RECT 141.930 57.600 142.190 57.650 ;
        RECT 142.840 57.600 143.240 57.650 ;
        RECT 144.755 57.600 145.015 57.650 ;
        RECT 145.280 57.600 145.540 57.650 ;
        RECT 4.620 56.585 5.000 56.985 ;
        RECT 16.590 56.600 17.060 56.970 ;
        RECT 22.775 56.925 23.100 57.105 ;
        RECT 139.740 56.950 140.040 57.500 ;
        RECT 148.740 57.410 149.840 58.490 ;
        RECT 151.540 57.625 151.975 58.475 ;
        RECT 155.255 56.975 155.420 194.030 ;
        RECT 24.075 56.925 24.425 56.950 ;
        RECT 22.775 56.605 24.465 56.925 ;
        RECT 24.035 56.580 24.465 56.605 ;
        RECT 139.690 56.600 140.090 56.950 ;
        RECT 146.320 56.580 146.760 56.970 ;
        RECT 155.040 56.575 155.420 56.975 ;
        RECT 25.295 55.060 26.345 55.110 ;
        RECT 25.295 54.060 26.350 55.060 ;
        RECT 133.640 55.000 134.640 56.000 ;
        RECT 25.295 54.010 26.345 54.060 ;
        RECT 8.850 51.710 24.185 53.210 ;
        RECT 25.295 53.060 26.345 53.110 ;
        RECT 25.295 52.060 26.350 53.060 ;
        RECT 25.295 52.010 26.345 52.060 ;
        RECT 133.640 51.700 147.725 53.200 ;
        RECT 25.300 51.010 26.350 51.060 ;
        RECT 11.950 49.510 26.350 51.010 ;
        RECT 8.065 47.635 8.500 48.485 ;
        RECT 10.200 47.420 11.245 48.500 ;
        RECT 16.815 48.010 17.235 48.460 ;
        RECT 17.865 48.010 18.125 48.060 ;
        RECT 18.390 48.010 18.650 48.060 ;
        RECT 19.300 48.010 19.700 48.060 ;
        RECT 21.215 48.010 21.475 48.060 ;
        RECT 21.740 48.010 22.000 48.060 ;
        RECT 22.670 48.010 23.200 48.060 ;
        RECT 24.640 48.010 24.940 49.510 ;
        RECT 25.300 49.460 26.350 49.510 ;
        RECT 133.640 49.400 134.690 50.500 ;
        RECT 135.490 49.500 151.190 51.000 ;
        RECT 134.390 49.000 134.690 49.400 ;
        RECT 134.390 48.700 135.540 49.000 ;
        RECT 16.815 47.660 18.125 48.010 ;
        RECT 18.350 47.660 21.500 48.010 ;
        RECT 21.725 47.660 24.125 48.010 ;
        RECT 24.390 47.660 24.940 48.010 ;
        RECT 17.865 47.610 18.125 47.660 ;
        RECT 18.390 47.610 18.650 47.660 ;
        RECT 19.300 47.610 19.700 47.660 ;
        RECT 21.215 47.425 21.475 47.660 ;
        RECT 21.740 47.610 22.000 47.660 ;
        RECT 21.215 47.105 23.100 47.425 ;
        RECT 25.200 47.420 26.350 48.500 ;
        RECT 133.640 47.400 134.690 48.500 ;
        RECT 135.240 47.800 135.540 48.700 ;
        RECT 140.355 48.000 140.775 48.450 ;
        RECT 141.405 48.000 141.665 48.050 ;
        RECT 141.930 48.000 142.190 48.050 ;
        RECT 142.840 48.000 143.240 48.050 ;
        RECT 144.755 48.000 145.015 48.050 ;
        RECT 145.280 48.000 145.540 48.050 ;
        RECT 146.840 48.000 147.340 48.460 ;
        RECT 135.240 47.500 140.040 47.800 ;
        RECT 140.355 47.650 141.665 48.000 ;
        RECT 141.890 47.650 145.040 48.000 ;
        RECT 145.265 47.650 147.340 48.000 ;
        RECT 141.405 47.600 141.665 47.650 ;
        RECT 141.930 47.600 142.190 47.650 ;
        RECT 142.840 47.600 143.240 47.650 ;
        RECT 144.755 47.600 145.015 47.650 ;
        RECT 145.280 47.600 145.540 47.650 ;
        RECT 4.295 46.585 4.675 46.985 ;
        RECT 16.590 46.600 17.060 46.970 ;
        RECT 22.775 46.925 23.100 47.105 ;
        RECT 139.740 46.950 140.040 47.500 ;
        RECT 148.740 47.410 149.840 48.490 ;
        RECT 151.540 47.625 151.975 48.475 ;
        RECT 155.580 46.975 155.745 194.690 ;
        RECT 24.075 46.925 24.425 46.950 ;
        RECT 22.775 46.605 24.465 46.925 ;
        RECT 24.035 46.580 24.465 46.605 ;
        RECT 139.690 46.600 140.090 46.950 ;
        RECT 146.320 46.580 146.760 46.970 ;
        RECT 155.365 46.575 155.745 46.975 ;
        RECT 25.295 45.060 26.345 45.110 ;
        RECT 25.295 44.060 26.350 45.060 ;
        RECT 133.640 45.000 134.640 46.000 ;
        RECT 25.295 44.010 26.345 44.060 ;
        RECT 8.850 41.710 24.185 43.210 ;
        RECT 25.295 43.060 26.345 43.110 ;
        RECT 25.295 42.060 26.350 43.060 ;
        RECT 25.295 42.010 26.345 42.060 ;
        RECT 133.640 41.700 147.725 43.200 ;
        RECT 25.300 41.010 26.350 41.060 ;
        RECT 11.950 39.510 26.350 41.010 ;
        RECT 8.065 37.635 8.500 38.485 ;
        RECT 10.200 37.420 11.245 38.500 ;
        RECT 16.815 38.010 17.235 38.460 ;
        RECT 17.865 38.010 18.125 38.060 ;
        RECT 18.390 38.010 18.650 38.060 ;
        RECT 19.300 38.010 19.700 38.060 ;
        RECT 21.215 38.010 21.475 38.060 ;
        RECT 21.740 38.010 22.000 38.060 ;
        RECT 22.670 38.010 23.200 38.060 ;
        RECT 24.640 38.010 24.940 39.510 ;
        RECT 25.300 39.460 26.350 39.510 ;
        RECT 133.640 39.400 134.690 40.500 ;
        RECT 135.490 39.500 151.190 41.000 ;
        RECT 134.390 39.000 134.690 39.400 ;
        RECT 134.390 38.700 135.540 39.000 ;
        RECT 16.815 37.660 18.125 38.010 ;
        RECT 18.350 37.660 21.500 38.010 ;
        RECT 21.725 37.660 24.125 38.010 ;
        RECT 24.390 37.660 24.940 38.010 ;
        RECT 17.865 37.610 18.125 37.660 ;
        RECT 18.390 37.610 18.650 37.660 ;
        RECT 19.300 37.610 19.700 37.660 ;
        RECT 21.215 37.425 21.475 37.660 ;
        RECT 21.740 37.610 22.000 37.660 ;
        RECT 21.215 37.105 23.100 37.425 ;
        RECT 25.200 37.420 26.350 38.500 ;
        RECT 133.640 37.400 134.690 38.500 ;
        RECT 135.240 37.800 135.540 38.700 ;
        RECT 140.355 38.000 140.775 38.450 ;
        RECT 141.405 38.000 141.665 38.050 ;
        RECT 141.930 38.000 142.190 38.050 ;
        RECT 142.840 38.000 143.240 38.050 ;
        RECT 144.755 38.000 145.015 38.050 ;
        RECT 145.280 38.000 145.540 38.050 ;
        RECT 146.840 38.000 147.340 38.460 ;
        RECT 135.240 37.500 140.040 37.800 ;
        RECT 140.355 37.650 141.665 38.000 ;
        RECT 141.890 37.650 145.040 38.000 ;
        RECT 145.265 37.650 147.340 38.000 ;
        RECT 141.405 37.600 141.665 37.650 ;
        RECT 141.930 37.600 142.190 37.650 ;
        RECT 142.840 37.600 143.240 37.650 ;
        RECT 144.755 37.600 145.015 37.650 ;
        RECT 145.280 37.600 145.540 37.650 ;
        RECT 3.970 36.585 4.350 36.985 ;
        RECT 16.590 36.600 17.060 36.970 ;
        RECT 22.775 36.925 23.100 37.105 ;
        RECT 139.740 36.950 140.040 37.500 ;
        RECT 148.740 37.410 149.840 38.490 ;
        RECT 151.540 37.625 151.975 38.475 ;
        RECT 155.905 36.975 156.070 195.350 ;
        RECT 24.075 36.925 24.425 36.950 ;
        RECT 22.775 36.605 24.465 36.925 ;
        RECT 24.035 36.580 24.465 36.605 ;
        RECT 139.690 36.600 140.090 36.950 ;
        RECT 146.320 36.580 146.760 36.970 ;
        RECT 155.690 36.575 156.070 36.975 ;
        RECT 25.295 35.060 26.345 35.110 ;
        RECT 25.295 34.060 26.350 35.060 ;
        RECT 133.640 35.000 134.640 36.000 ;
        RECT 25.295 34.010 26.345 34.060 ;
        RECT 8.850 31.710 24.185 33.210 ;
        RECT 25.295 33.060 26.345 33.110 ;
        RECT 25.295 32.060 26.350 33.060 ;
        RECT 25.295 32.010 26.345 32.060 ;
        RECT 133.640 31.700 147.725 33.200 ;
        RECT 25.300 31.010 26.350 31.060 ;
        RECT 11.950 29.510 26.350 31.010 ;
        RECT 8.065 27.635 8.500 28.485 ;
        RECT 10.200 27.420 11.245 28.500 ;
        RECT 16.815 28.010 17.235 28.460 ;
        RECT 17.865 28.010 18.125 28.060 ;
        RECT 18.390 28.010 18.650 28.060 ;
        RECT 19.300 28.010 19.700 28.060 ;
        RECT 21.215 28.010 21.475 28.060 ;
        RECT 21.740 28.010 22.000 28.060 ;
        RECT 22.670 28.010 23.200 28.060 ;
        RECT 24.640 28.010 24.940 29.510 ;
        RECT 25.300 29.460 26.350 29.510 ;
        RECT 133.640 29.400 134.690 30.500 ;
        RECT 135.490 29.500 151.190 31.000 ;
        RECT 134.390 29.000 134.690 29.400 ;
        RECT 134.390 28.700 135.540 29.000 ;
        RECT 16.815 27.660 18.125 28.010 ;
        RECT 18.350 27.660 21.500 28.010 ;
        RECT 21.725 27.660 24.125 28.010 ;
        RECT 24.390 27.660 24.940 28.010 ;
        RECT 17.865 27.610 18.125 27.660 ;
        RECT 18.390 27.610 18.650 27.660 ;
        RECT 19.300 27.610 19.700 27.660 ;
        RECT 21.215 27.425 21.475 27.660 ;
        RECT 21.740 27.610 22.000 27.660 ;
        RECT 21.215 27.105 23.100 27.425 ;
        RECT 25.200 27.420 26.350 28.500 ;
        RECT 133.640 27.400 134.690 28.500 ;
        RECT 135.240 27.800 135.540 28.700 ;
        RECT 140.355 28.000 140.775 28.450 ;
        RECT 141.405 28.000 141.665 28.050 ;
        RECT 141.930 28.000 142.190 28.050 ;
        RECT 142.840 28.000 143.240 28.050 ;
        RECT 144.755 28.000 145.015 28.050 ;
        RECT 145.280 28.000 145.540 28.050 ;
        RECT 146.840 28.000 147.340 28.460 ;
        RECT 135.240 27.500 140.040 27.800 ;
        RECT 140.355 27.650 141.665 28.000 ;
        RECT 141.890 27.650 145.040 28.000 ;
        RECT 145.265 27.650 147.340 28.000 ;
        RECT 141.405 27.600 141.665 27.650 ;
        RECT 141.930 27.600 142.190 27.650 ;
        RECT 142.840 27.600 143.240 27.650 ;
        RECT 144.755 27.600 145.015 27.650 ;
        RECT 145.280 27.600 145.540 27.650 ;
        RECT 3.645 26.585 4.025 26.985 ;
        RECT 16.590 26.600 17.060 26.970 ;
        RECT 22.775 26.925 23.100 27.105 ;
        RECT 139.740 26.950 140.040 27.500 ;
        RECT 148.740 27.410 149.840 28.490 ;
        RECT 151.540 27.625 151.975 28.475 ;
        RECT 156.230 26.975 156.395 196.010 ;
        RECT 24.075 26.925 24.425 26.950 ;
        RECT 22.775 26.605 24.465 26.925 ;
        RECT 24.035 26.580 24.465 26.605 ;
        RECT 139.690 26.600 140.090 26.950 ;
        RECT 146.320 26.580 146.760 26.970 ;
        RECT 156.015 26.575 156.395 26.975 ;
        RECT 25.295 25.060 26.345 25.110 ;
        RECT 25.295 24.060 26.350 25.060 ;
        RECT 133.640 25.000 134.640 26.000 ;
        RECT 25.295 24.010 26.345 24.060 ;
        RECT 8.850 21.710 24.185 23.210 ;
        RECT 25.295 23.060 26.345 23.110 ;
        RECT 25.295 22.060 26.350 23.060 ;
        RECT 25.295 22.010 26.345 22.060 ;
        RECT 133.640 21.700 147.725 23.200 ;
        RECT 25.300 21.010 26.350 21.060 ;
        RECT 11.950 19.510 26.350 21.010 ;
        RECT 8.065 17.635 8.500 18.485 ;
        RECT 10.200 17.420 11.245 18.500 ;
        RECT 16.815 18.010 17.235 18.460 ;
        RECT 17.865 18.010 18.125 18.060 ;
        RECT 18.390 18.010 18.650 18.060 ;
        RECT 19.300 18.010 19.700 18.060 ;
        RECT 21.215 18.010 21.475 18.060 ;
        RECT 21.740 18.010 22.000 18.060 ;
        RECT 22.670 18.010 23.200 18.060 ;
        RECT 24.640 18.010 24.940 19.510 ;
        RECT 25.300 19.460 26.350 19.510 ;
        RECT 133.640 19.400 134.690 20.500 ;
        RECT 135.490 19.500 151.190 21.000 ;
        RECT 134.390 19.000 134.690 19.400 ;
        RECT 134.390 18.700 135.540 19.000 ;
        RECT 16.815 17.660 18.125 18.010 ;
        RECT 18.350 17.660 21.500 18.010 ;
        RECT 21.725 17.660 24.125 18.010 ;
        RECT 24.390 17.660 24.940 18.010 ;
        RECT 17.865 17.610 18.125 17.660 ;
        RECT 18.390 17.610 18.650 17.660 ;
        RECT 19.300 17.610 19.700 17.660 ;
        RECT 21.215 17.425 21.475 17.660 ;
        RECT 21.740 17.610 22.000 17.660 ;
        RECT 21.215 17.105 23.100 17.425 ;
        RECT 25.200 17.420 26.350 18.500 ;
        RECT 133.640 17.400 134.690 18.500 ;
        RECT 135.240 17.800 135.540 18.700 ;
        RECT 140.355 18.000 140.775 18.450 ;
        RECT 141.405 18.000 141.665 18.050 ;
        RECT 141.930 18.000 142.190 18.050 ;
        RECT 142.840 18.000 143.240 18.050 ;
        RECT 144.755 18.000 145.015 18.050 ;
        RECT 145.280 18.000 145.540 18.050 ;
        RECT 146.840 18.000 147.340 18.460 ;
        RECT 135.240 17.500 140.040 17.800 ;
        RECT 140.355 17.650 141.665 18.000 ;
        RECT 141.890 17.650 145.040 18.000 ;
        RECT 145.265 17.650 147.340 18.000 ;
        RECT 141.405 17.600 141.665 17.650 ;
        RECT 141.930 17.600 142.190 17.650 ;
        RECT 142.840 17.600 143.240 17.650 ;
        RECT 144.755 17.600 145.015 17.650 ;
        RECT 145.280 17.600 145.540 17.650 ;
        RECT 3.320 16.585 3.700 16.985 ;
        RECT 16.590 16.600 17.060 16.970 ;
        RECT 22.775 16.925 23.100 17.105 ;
        RECT 139.740 16.950 140.040 17.500 ;
        RECT 148.740 17.410 149.840 18.490 ;
        RECT 151.540 17.625 151.975 18.475 ;
        RECT 156.555 16.975 156.720 196.670 ;
        RECT 24.075 16.925 24.425 16.950 ;
        RECT 22.775 16.605 24.465 16.925 ;
        RECT 24.035 16.580 24.465 16.605 ;
        RECT 139.690 16.600 140.090 16.950 ;
        RECT 146.320 16.580 146.760 16.970 ;
        RECT 156.340 16.575 156.720 16.975 ;
        RECT 25.295 15.060 26.345 15.110 ;
        RECT 25.295 14.060 26.350 15.060 ;
        RECT 133.640 15.000 134.640 16.000 ;
        RECT 25.295 14.010 26.345 14.060 ;
        RECT 8.850 11.710 24.185 13.210 ;
        RECT 25.295 13.060 26.345 13.110 ;
        RECT 25.295 12.060 26.350 13.060 ;
        RECT 25.295 12.010 26.345 12.060 ;
        RECT 133.640 11.700 147.725 13.200 ;
        RECT 25.300 11.010 26.350 11.060 ;
        RECT 11.950 9.510 26.350 11.010 ;
        RECT 8.065 7.635 8.500 8.485 ;
        RECT 10.200 7.420 11.245 8.500 ;
        RECT 16.815 8.010 17.235 8.460 ;
        RECT 17.865 8.010 18.125 8.060 ;
        RECT 18.390 8.010 18.650 8.060 ;
        RECT 19.300 8.010 19.700 8.060 ;
        RECT 21.215 8.010 21.475 8.060 ;
        RECT 21.740 8.010 22.000 8.060 ;
        RECT 22.670 8.010 23.200 8.060 ;
        RECT 24.640 8.010 24.940 9.510 ;
        RECT 25.300 9.460 26.350 9.510 ;
        RECT 133.640 9.400 134.690 10.500 ;
        RECT 135.490 9.500 151.190 11.000 ;
        RECT 134.390 9.000 134.690 9.400 ;
        RECT 134.390 8.700 135.540 9.000 ;
        RECT 16.815 7.660 18.125 8.010 ;
        RECT 18.350 7.660 21.500 8.010 ;
        RECT 21.725 7.660 24.125 8.010 ;
        RECT 24.390 7.660 24.940 8.010 ;
        RECT 17.865 7.610 18.125 7.660 ;
        RECT 18.390 7.610 18.650 7.660 ;
        RECT 19.300 7.610 19.700 7.660 ;
        RECT 21.215 7.425 21.475 7.660 ;
        RECT 21.740 7.610 22.000 7.660 ;
        RECT 21.215 7.105 23.100 7.425 ;
        RECT 25.200 7.420 26.350 8.500 ;
        RECT 133.640 7.400 134.690 8.500 ;
        RECT 135.240 7.800 135.540 8.700 ;
        RECT 140.355 8.000 140.775 8.450 ;
        RECT 141.405 8.000 141.665 8.050 ;
        RECT 141.930 8.000 142.190 8.050 ;
        RECT 142.840 8.000 143.240 8.050 ;
        RECT 144.755 8.000 145.015 8.050 ;
        RECT 145.280 8.000 145.540 8.050 ;
        RECT 146.840 8.000 147.340 8.460 ;
        RECT 135.240 7.500 140.040 7.800 ;
        RECT 140.355 7.650 141.665 8.000 ;
        RECT 141.890 7.650 145.040 8.000 ;
        RECT 145.265 7.650 147.340 8.000 ;
        RECT 141.405 7.600 141.665 7.650 ;
        RECT 141.930 7.600 142.190 7.650 ;
        RECT 142.840 7.600 143.240 7.650 ;
        RECT 144.755 7.600 145.015 7.650 ;
        RECT 145.280 7.600 145.540 7.650 ;
        RECT 2.995 6.585 3.375 6.985 ;
        RECT 16.590 6.600 17.060 6.970 ;
        RECT 22.775 6.925 23.100 7.105 ;
        RECT 139.740 6.950 140.040 7.500 ;
        RECT 148.740 7.410 149.840 8.490 ;
        RECT 151.540 7.625 151.975 8.475 ;
        RECT 156.880 6.975 157.045 197.330 ;
        RECT 24.075 6.925 24.425 6.950 ;
        RECT 22.775 6.605 24.465 6.925 ;
        RECT 24.035 6.580 24.465 6.605 ;
        RECT 139.690 6.600 140.090 6.950 ;
        RECT 146.320 6.580 146.760 6.970 ;
        RECT 156.665 6.575 157.045 6.975 ;
        RECT 157.205 5.990 157.370 197.990 ;
        RECT 157.570 197.410 158.880 198.820 ;
      LAYER met3 ;
        RECT 22.605 224.130 22.935 224.135 ;
        RECT 22.350 224.120 22.935 224.130 ;
        RECT 79.185 224.120 79.515 224.135 ;
        RECT 81.230 224.120 81.610 224.130 ;
        RECT 22.350 223.820 23.160 224.120 ;
        RECT 79.185 223.820 81.610 224.120 ;
        RECT 22.350 223.810 22.935 223.820 ;
        RECT 22.605 223.805 22.935 223.810 ;
        RECT 79.185 223.805 79.515 223.820 ;
        RECT 81.230 223.810 81.610 223.820 ;
        RECT 85.165 224.120 85.495 224.135 ;
        RECT 88.590 224.120 88.970 224.130 ;
        RECT 85.165 223.820 88.970 224.120 ;
        RECT 85.165 223.805 85.495 223.820 ;
        RECT 88.590 223.810 88.970 223.820 ;
        RECT 121.710 224.120 122.090 224.130 ;
        RECT 126.105 224.120 126.435 224.135 ;
        RECT 121.710 223.820 126.435 224.120 ;
        RECT 121.710 223.810 122.090 223.820 ;
        RECT 126.105 223.805 126.435 223.820 ;
        RECT 48.365 223.450 48.695 223.455 ;
        RECT 48.110 223.440 48.695 223.450 ;
        RECT 40.840 222.875 42.420 223.205 ;
        RECT 47.910 223.140 48.695 223.440 ;
        RECT 125.390 223.440 125.770 223.450 ;
        RECT 127.485 223.440 127.815 223.455 ;
        RECT 48.110 223.130 48.695 223.140 ;
        RECT 48.365 223.125 48.695 223.130 ;
        RECT 79.710 222.875 81.290 223.205 ;
        RECT 118.580 222.875 120.160 223.205 ;
        RECT 125.390 223.140 127.815 223.440 ;
        RECT 125.390 223.130 125.770 223.140 ;
        RECT 127.485 223.125 127.815 223.140 ;
        RECT 132.750 223.440 133.130 223.450 ;
        RECT 133.925 223.440 134.255 223.455 ;
        RECT 132.750 223.140 134.255 223.440 ;
        RECT 132.750 223.130 133.130 223.140 ;
        RECT 133.925 223.125 134.255 223.140 ;
        RECT 136.430 223.440 136.810 223.450 ;
        RECT 143.125 223.440 143.455 223.455 ;
        RECT 136.430 223.140 143.455 223.440 ;
        RECT 136.430 223.130 136.810 223.140 ;
        RECT 143.125 223.125 143.455 223.140 ;
        RECT 157.450 222.875 159.030 223.205 ;
        RECT 4.205 222.770 4.535 222.775 ;
        RECT 7.885 222.770 8.215 222.775 ;
        RECT 11.565 222.770 11.895 222.775 ;
        RECT 3.950 222.760 4.535 222.770 ;
        RECT 7.630 222.760 8.215 222.770 ;
        RECT 11.310 222.760 11.895 222.770 ;
        RECT 14.990 222.760 15.370 222.770 ;
        RECT 16.165 222.760 16.495 222.775 ;
        RECT 18.925 222.770 19.255 222.775 ;
        RECT 26.285 222.770 26.615 222.775 ;
        RECT 29.965 222.770 30.295 222.775 ;
        RECT 3.950 222.460 4.760 222.760 ;
        RECT 7.630 222.460 8.440 222.760 ;
        RECT 11.310 222.460 12.120 222.760 ;
        RECT 14.990 222.460 16.495 222.760 ;
        RECT 3.950 222.450 4.535 222.460 ;
        RECT 7.630 222.450 8.215 222.460 ;
        RECT 11.310 222.450 11.895 222.460 ;
        RECT 14.990 222.450 15.370 222.460 ;
        RECT 4.205 222.445 4.535 222.450 ;
        RECT 7.885 222.445 8.215 222.450 ;
        RECT 11.565 222.445 11.895 222.450 ;
        RECT 16.165 222.445 16.495 222.460 ;
        RECT 18.670 222.760 19.255 222.770 ;
        RECT 26.030 222.760 26.615 222.770 ;
        RECT 29.710 222.760 30.295 222.770 ;
        RECT 62.830 222.760 63.210 222.770 ;
        RECT 70.445 222.760 70.775 222.775 ;
        RECT 18.670 222.460 19.480 222.760 ;
        RECT 26.030 222.460 26.840 222.760 ;
        RECT 29.710 222.460 30.520 222.760 ;
        RECT 62.830 222.460 70.775 222.760 ;
        RECT 18.670 222.450 19.255 222.460 ;
        RECT 26.030 222.450 26.615 222.460 ;
        RECT 29.710 222.450 30.295 222.460 ;
        RECT 62.830 222.450 63.210 222.460 ;
        RECT 18.925 222.445 19.255 222.450 ;
        RECT 26.285 222.445 26.615 222.450 ;
        RECT 29.965 222.445 30.295 222.450 ;
        RECT 70.445 222.445 70.775 222.460 ;
        RECT 73.665 222.080 73.995 222.095 ;
        RECT 77.550 222.080 77.930 222.090 ;
        RECT 73.665 221.780 77.930 222.080 ;
        RECT 73.665 221.765 73.995 221.780 ;
        RECT 77.550 221.770 77.930 221.780 ;
        RECT 84.910 222.080 85.290 222.090 ;
        RECT 87.005 222.080 87.335 222.095 ;
        RECT 84.910 221.780 87.335 222.080 ;
        RECT 84.910 221.770 85.290 221.780 ;
        RECT 87.005 221.765 87.335 221.780 ;
        RECT 140.365 220.730 140.695 220.735 ;
        RECT 147.725 220.730 148.055 220.735 ;
        RECT 140.110 220.720 140.695 220.730 ;
        RECT 147.470 220.720 148.055 220.730 ;
        RECT 1.010 220.155 2.590 220.485 ;
        RECT 21.405 220.155 22.985 220.485 ;
        RECT 60.275 220.155 61.855 220.485 ;
        RECT 99.145 220.155 100.725 220.485 ;
        RECT 138.015 220.155 139.595 220.485 ;
        RECT 140.110 220.420 140.920 220.720 ;
        RECT 147.270 220.420 148.055 220.720 ;
        RECT 140.110 220.410 140.695 220.420 ;
        RECT 147.470 220.410 148.055 220.420 ;
        RECT 140.365 220.405 140.695 220.410 ;
        RECT 147.725 220.405 148.055 220.410 ;
        RECT 108.625 220.040 108.955 220.055 ;
        RECT 118.285 220.040 118.615 220.055 ;
        RECT 108.625 219.740 118.615 220.040 ;
        RECT 108.625 219.725 108.955 219.740 ;
        RECT 118.285 219.725 118.615 219.740 ;
        RECT 154.625 220.050 154.955 220.055 ;
        RECT 154.625 220.040 155.210 220.050 ;
        RECT 154.625 219.740 155.410 220.040 ;
        RECT 154.625 219.730 155.210 219.740 ;
        RECT 154.625 219.725 154.955 219.730 ;
        RECT 69.985 219.370 70.315 219.375 ;
        RECT 144.045 219.370 144.375 219.375 ;
        RECT 69.985 219.360 70.570 219.370 ;
        RECT 143.790 219.360 144.375 219.370 ;
        RECT 69.760 219.060 70.570 219.360 ;
        RECT 143.590 219.060 144.375 219.360 ;
        RECT 69.985 219.050 70.570 219.060 ;
        RECT 143.790 219.050 144.375 219.060 ;
        RECT 69.985 219.045 70.315 219.050 ;
        RECT 144.045 219.045 144.375 219.050 ;
        RECT 40.840 217.435 42.420 217.765 ;
        RECT 79.710 217.435 81.290 217.765 ;
        RECT 118.580 217.435 120.160 217.765 ;
        RECT 157.450 217.435 159.030 217.765 ;
        RECT 70.905 216.640 71.235 216.655 ;
        RECT 73.870 216.640 74.250 216.650 ;
        RECT 70.905 216.340 74.250 216.640 ;
        RECT 70.905 216.325 71.235 216.340 ;
        RECT 73.870 216.330 74.250 216.340 ;
        RECT 74.585 216.640 74.915 216.655 ;
        RECT 85.625 216.640 85.955 216.655 ;
        RECT 74.585 216.340 85.955 216.640 ;
        RECT 74.585 216.325 74.915 216.340 ;
        RECT 85.625 216.325 85.955 216.340 ;
        RECT 99.425 215.960 99.755 215.975 ;
        RECT 112.305 215.960 112.635 215.975 ;
        RECT 126.105 215.960 126.435 215.975 ;
        RECT 130.245 215.960 130.575 215.975 ;
        RECT 99.425 215.660 130.575 215.960 ;
        RECT 99.425 215.645 99.755 215.660 ;
        RECT 112.305 215.645 112.635 215.660 ;
        RECT 126.105 215.645 126.435 215.660 ;
        RECT 130.245 215.645 130.575 215.660 ;
        RECT 1.010 214.715 2.590 215.045 ;
        RECT 21.405 214.715 22.985 215.045 ;
        RECT 60.275 214.715 61.855 215.045 ;
        RECT 99.145 214.715 100.725 215.045 ;
        RECT 138.015 214.715 139.595 215.045 ;
        RECT 55.725 213.920 56.055 213.935 ;
        RECT 85.165 213.920 85.495 213.935 ;
        RECT 55.725 213.620 85.495 213.920 ;
        RECT 55.725 213.605 56.055 213.620 ;
        RECT 85.165 213.605 85.495 213.620 ;
        RECT 59.865 213.240 60.195 213.255 ;
        RECT 64.925 213.240 65.255 213.255 ;
        RECT 59.865 212.940 65.255 213.240 ;
        RECT 59.865 212.925 60.195 212.940 ;
        RECT 64.925 212.925 65.255 212.940 ;
        RECT 71.825 213.240 72.155 213.255 ;
        RECT 78.725 213.240 79.055 213.255 ;
        RECT 91.145 213.240 91.475 213.255 ;
        RECT 71.825 212.940 91.475 213.240 ;
        RECT 71.825 212.925 72.155 212.940 ;
        RECT 78.725 212.925 79.055 212.940 ;
        RECT 91.145 212.925 91.475 212.940 ;
        RECT 40.840 211.995 42.420 212.325 ;
        RECT 79.710 211.995 81.290 212.325 ;
        RECT 118.580 211.995 120.160 212.325 ;
        RECT 157.450 211.995 159.030 212.325 ;
        RECT 62.165 211.880 62.495 211.895 ;
        RECT 66.510 211.880 66.890 211.890 ;
        RECT 62.165 211.580 66.890 211.880 ;
        RECT 62.165 211.565 62.495 211.580 ;
        RECT 66.510 211.570 66.890 211.580 ;
        RECT 37.070 211.200 37.450 211.210 ;
        RECT 55.725 211.200 56.055 211.215 ;
        RECT 86.085 211.200 86.415 211.215 ;
        RECT 37.070 210.900 56.055 211.200 ;
        RECT 37.070 210.890 37.450 210.900 ;
        RECT 55.725 210.885 56.055 210.900 ;
        RECT 56.430 210.900 86.415 211.200 ;
        RECT 56.430 210.535 56.730 210.900 ;
        RECT 86.085 210.885 86.415 210.900 ;
        RECT 98.965 211.200 99.295 211.215 ;
        RECT 101.265 211.200 101.595 211.215 ;
        RECT 104.945 211.200 105.275 211.215 ;
        RECT 98.965 210.900 105.275 211.200 ;
        RECT 98.965 210.885 99.295 210.900 ;
        RECT 101.265 210.885 101.595 210.900 ;
        RECT 104.945 210.885 105.275 210.900 ;
        RECT 113.225 211.200 113.555 211.215 ;
        RECT 151.150 211.200 151.530 211.210 ;
        RECT 113.225 210.900 151.530 211.200 ;
        RECT 113.225 210.885 113.555 210.900 ;
        RECT 151.150 210.890 151.530 210.900 ;
        RECT 39.830 210.520 40.210 210.530 ;
        RECT 56.185 210.520 56.730 210.535 ;
        RECT 77.805 210.520 78.135 210.535 ;
        RECT 39.830 210.220 56.730 210.520 ;
        RECT 57.350 210.220 78.135 210.520 ;
        RECT 39.830 210.210 40.210 210.220 ;
        RECT 56.185 210.205 56.515 210.220 ;
        RECT 51.790 209.840 52.170 209.850 ;
        RECT 57.350 209.840 57.650 210.220 ;
        RECT 77.805 210.205 78.135 210.220 ;
        RECT 81.025 210.520 81.355 210.535 ;
        RECT 85.625 210.520 85.955 210.535 ;
        RECT 81.025 210.220 85.955 210.520 ;
        RECT 81.025 210.205 81.355 210.220 ;
        RECT 85.625 210.205 85.955 210.220 ;
        RECT 97.125 210.520 97.455 210.535 ;
        RECT 104.025 210.520 104.355 210.535 ;
        RECT 97.125 210.220 104.355 210.520 ;
        RECT 97.125 210.205 97.455 210.220 ;
        RECT 104.025 210.205 104.355 210.220 ;
        RECT 1.010 209.275 2.590 209.605 ;
        RECT 21.405 209.275 22.985 209.605 ;
        RECT 51.790 209.540 57.650 209.840 ;
        RECT 75.505 209.840 75.835 209.855 ;
        RECT 87.005 209.840 87.335 209.855 ;
        RECT 51.790 209.530 52.170 209.540 ;
        RECT 60.275 209.275 61.855 209.605 ;
        RECT 75.505 209.540 87.335 209.840 ;
        RECT 75.505 209.525 75.835 209.540 ;
        RECT 87.005 209.525 87.335 209.540 ;
        RECT 99.145 209.275 100.725 209.605 ;
        RECT 138.015 209.275 139.595 209.605 ;
        RECT 44.430 209.160 44.810 209.170 ;
        RECT 59.405 209.160 59.735 209.175 ;
        RECT 44.430 208.860 59.735 209.160 ;
        RECT 44.430 208.850 44.810 208.860 ;
        RECT 59.405 208.845 59.735 208.860 ;
        RECT 75.965 209.160 76.295 209.175 ;
        RECT 82.405 209.160 82.735 209.175 ;
        RECT 75.965 208.860 82.735 209.160 ;
        RECT 75.965 208.845 76.295 208.860 ;
        RECT 82.405 208.845 82.735 208.860 ;
        RECT 153.705 209.160 154.035 209.175 ;
        RECT 156.670 209.160 157.050 209.170 ;
        RECT 153.705 208.860 157.050 209.160 ;
        RECT 153.705 208.845 154.035 208.860 ;
        RECT 156.670 208.850 157.050 208.860 ;
        RECT 33.390 208.480 33.770 208.490 ;
        RECT 65.385 208.480 65.715 208.495 ;
        RECT 33.390 208.180 65.715 208.480 ;
        RECT 33.390 208.170 33.770 208.180 ;
        RECT 65.385 208.165 65.715 208.180 ;
        RECT 66.305 208.480 66.635 208.495 ;
        RECT 101.725 208.480 102.055 208.495 ;
        RECT 66.305 208.180 102.055 208.480 ;
        RECT 66.305 208.165 66.635 208.180 ;
        RECT 101.725 208.165 102.055 208.180 ;
        RECT 23.270 207.800 23.650 207.810 ;
        RECT 62.625 207.800 62.955 207.815 ;
        RECT 23.270 207.500 62.955 207.800 ;
        RECT 23.270 207.490 23.650 207.500 ;
        RECT 62.625 207.485 62.955 207.500 ;
        RECT 64.925 207.800 65.255 207.815 ;
        RECT 69.985 207.800 70.315 207.815 ;
        RECT 87.465 207.800 87.795 207.815 ;
        RECT 107.245 207.800 107.575 207.815 ;
        RECT 64.925 207.500 70.315 207.800 ;
        RECT 64.925 207.485 65.255 207.500 ;
        RECT 69.985 207.485 70.315 207.500 ;
        RECT 78.740 207.500 107.575 207.800 ;
        RECT 55.470 207.120 55.850 207.130 ;
        RECT 78.740 207.120 79.040 207.500 ;
        RECT 87.465 207.485 87.795 207.500 ;
        RECT 107.245 207.485 107.575 207.500 ;
        RECT 40.840 206.555 42.420 206.885 ;
        RECT 55.470 206.820 79.040 207.120 ;
        RECT 84.245 207.120 84.575 207.135 ;
        RECT 86.545 207.120 86.875 207.135 ;
        RECT 55.470 206.810 55.850 206.820 ;
        RECT 79.710 206.555 81.290 206.885 ;
        RECT 84.245 206.820 86.875 207.120 ;
        RECT 84.245 206.805 84.575 206.820 ;
        RECT 86.545 206.805 86.875 206.820 ;
        RECT 118.580 206.555 120.160 206.885 ;
        RECT 157.450 206.555 159.030 206.885 ;
        RECT 48.110 206.440 48.490 206.450 ;
        RECT 58.485 206.440 58.815 206.455 ;
        RECT 48.110 206.140 58.815 206.440 ;
        RECT 48.110 206.130 48.490 206.140 ;
        RECT 58.485 206.125 58.815 206.140 ;
        RECT 59.150 206.440 59.530 206.450 ;
        RECT 59.150 206.140 79.040 206.440 ;
        RECT 59.150 206.130 59.530 206.140 ;
        RECT 6.710 205.760 7.090 205.770 ;
        RECT 10.645 205.760 10.975 205.775 ;
        RECT 6.710 205.460 10.975 205.760 ;
        RECT 6.710 205.450 7.090 205.460 ;
        RECT 10.645 205.445 10.975 205.460 ;
        RECT 14.070 205.760 14.450 205.770 ;
        RECT 21.685 205.760 22.015 205.775 ;
        RECT 14.070 205.460 22.015 205.760 ;
        RECT 14.070 205.450 14.450 205.460 ;
        RECT 21.685 205.445 22.015 205.460 ;
        RECT 28.790 205.760 29.170 205.770 ;
        RECT 32.725 205.760 33.055 205.775 ;
        RECT 28.790 205.460 33.055 205.760 ;
        RECT 28.790 205.450 29.170 205.460 ;
        RECT 32.725 205.445 33.055 205.460 ;
        RECT 36.150 205.760 36.530 205.770 ;
        RECT 40.085 205.760 40.415 205.775 ;
        RECT 36.150 205.460 40.415 205.760 ;
        RECT 36.150 205.450 36.530 205.460 ;
        RECT 40.085 205.445 40.415 205.460 ;
        RECT 55.470 205.760 55.850 205.770 ;
        RECT 58.945 205.760 59.275 205.775 ;
        RECT 55.470 205.460 59.275 205.760 ;
        RECT 55.470 205.450 55.850 205.460 ;
        RECT 58.945 205.445 59.275 205.460 ;
        RECT 63.085 205.760 63.415 205.775 ;
        RECT 71.365 205.760 71.695 205.775 ;
        RECT 77.805 205.770 78.135 205.775 ;
        RECT 77.550 205.760 78.135 205.770 ;
        RECT 63.085 205.460 71.695 205.760 ;
        RECT 77.350 205.460 78.135 205.760 ;
        RECT 78.740 205.760 79.040 206.140 ;
        RECT 80.565 205.760 80.895 205.775 ;
        RECT 88.385 205.760 88.715 205.775 ;
        RECT 78.740 205.460 88.715 205.760 ;
        RECT 63.085 205.445 63.415 205.460 ;
        RECT 71.365 205.445 71.695 205.460 ;
        RECT 77.550 205.450 78.135 205.460 ;
        RECT 77.805 205.445 78.135 205.450 ;
        RECT 80.565 205.445 80.895 205.460 ;
        RECT 88.385 205.445 88.715 205.460 ;
        RECT 89.765 205.760 90.095 205.775 ;
        RECT 92.270 205.760 92.650 205.770 ;
        RECT 89.765 205.460 92.650 205.760 ;
        RECT 89.765 205.445 90.095 205.460 ;
        RECT 92.270 205.450 92.650 205.460 ;
        RECT 103.105 205.760 103.435 205.775 ;
        RECT 114.145 205.770 114.475 205.775 ;
        RECT 106.990 205.760 107.370 205.770 ;
        RECT 103.105 205.460 107.370 205.760 ;
        RECT 103.105 205.445 103.435 205.460 ;
        RECT 106.990 205.450 107.370 205.460 ;
        RECT 114.145 205.760 114.730 205.770 ;
        RECT 117.825 205.760 118.155 205.775 ;
        RECT 128.865 205.770 129.195 205.775 ;
        RECT 150.945 205.770 151.275 205.775 ;
        RECT 121.710 205.760 122.090 205.770 ;
        RECT 114.145 205.460 114.930 205.760 ;
        RECT 117.825 205.460 122.090 205.760 ;
        RECT 114.145 205.450 114.730 205.460 ;
        RECT 114.145 205.445 114.475 205.450 ;
        RECT 117.825 205.445 118.155 205.460 ;
        RECT 121.710 205.450 122.090 205.460 ;
        RECT 128.865 205.760 129.450 205.770 ;
        RECT 150.945 205.760 151.530 205.770 ;
        RECT 128.865 205.460 129.650 205.760 ;
        RECT 150.945 205.460 151.730 205.760 ;
        RECT 128.865 205.450 129.450 205.460 ;
        RECT 150.945 205.450 151.530 205.460 ;
        RECT 128.865 205.445 129.195 205.450 ;
        RECT 150.945 205.445 151.275 205.450 ;
        RECT 1.010 203.835 2.590 204.165 ;
        RECT 21.405 203.835 22.985 204.165 ;
        RECT 60.275 203.835 61.855 204.165 ;
        RECT 99.145 203.835 100.725 204.165 ;
        RECT 138.015 203.835 139.595 204.165 ;
        RECT 136.225 201.690 136.555 201.695 ;
        RECT 136.225 201.680 136.810 201.690 ;
        RECT 40.840 201.115 42.420 201.445 ;
        RECT 79.710 201.115 81.290 201.445 ;
        RECT 118.580 201.115 120.160 201.445 ;
        RECT 136.225 201.380 137.010 201.680 ;
        RECT 136.225 201.370 136.810 201.380 ;
        RECT 136.225 201.365 136.555 201.370 ;
        RECT 157.450 201.115 159.030 201.445 ;
        RECT 70.190 201.000 70.570 201.010 ;
        RECT 71.825 201.000 72.155 201.015 ;
        RECT 70.190 200.700 72.155 201.000 ;
        RECT 70.190 200.690 70.570 200.700 ;
        RECT 71.825 200.685 72.155 200.700 ;
        RECT 143.585 201.010 143.915 201.015 ;
        RECT 143.585 201.000 144.170 201.010 ;
        RECT 143.585 200.700 144.370 201.000 ;
        RECT 143.585 200.690 144.170 200.700 ;
        RECT 143.585 200.685 143.915 200.690 ;
        RECT 62.830 200.320 63.210 200.330 ;
        RECT 64.005 200.320 64.335 200.335 ;
        RECT 40.640 199.810 42.610 200.270 ;
        RECT 62.830 200.020 64.335 200.320 ;
        RECT 62.830 200.010 63.210 200.020 ;
        RECT 64.005 200.005 64.335 200.020 ;
        RECT 84.705 200.330 85.035 200.335 ;
        RECT 84.705 200.320 85.290 200.330 ;
        RECT 84.705 200.020 85.490 200.320 ;
        RECT 84.705 200.010 85.290 200.020 ;
        RECT 84.705 200.005 85.035 200.010 ;
        RECT 5.250 198.980 5.790 199.010 ;
        RECT 6.880 198.980 7.270 199.015 ;
        RECT 5.250 198.680 7.270 198.980 ;
        RECT 5.250 198.630 5.790 198.680 ;
        RECT 6.880 198.625 7.270 198.680 ;
        RECT 14.240 199.010 14.630 199.020 ;
        RECT 14.240 198.630 15.400 199.010 ;
        RECT 14.240 198.625 14.630 198.630 ;
        RECT 2.670 198.320 3.030 198.350 ;
        RECT 151.145 198.320 151.525 198.370 ;
        RECT 157.010 198.320 157.370 198.350 ;
        RECT 2.670 198.020 157.370 198.320 ;
        RECT 2.670 197.990 3.030 198.020 ;
        RECT 157.010 197.990 157.370 198.020 ;
        RECT 2.995 197.660 3.355 197.690 ;
        RECT 143.785 197.660 144.165 197.710 ;
        RECT 156.685 197.660 157.045 197.690 ;
        RECT 2.995 197.360 157.050 197.660 ;
        RECT 157.670 197.410 158.880 198.820 ;
        RECT 2.995 197.330 3.355 197.360 ;
        RECT 156.685 197.330 157.045 197.360 ;
        RECT 3.320 197.000 3.680 197.030 ;
        RECT 136.425 197.000 136.805 197.050 ;
        RECT 156.360 197.000 156.720 197.030 ;
        RECT 3.320 196.700 156.725 197.000 ;
        RECT 3.320 196.670 3.680 196.700 ;
        RECT 156.360 196.670 156.720 196.700 ;
        RECT 3.645 196.340 4.005 196.370 ;
        RECT 129.065 196.340 129.445 196.390 ;
        RECT 156.035 196.340 156.395 196.370 ;
        RECT 3.645 196.040 156.400 196.340 ;
        RECT 3.645 196.010 4.005 196.040 ;
        RECT 156.035 196.010 156.395 196.040 ;
        RECT 3.970 195.680 4.330 195.710 ;
        RECT 121.705 195.680 122.085 195.730 ;
        RECT 155.710 195.680 156.070 195.710 ;
        RECT 3.970 195.380 156.075 195.680 ;
        RECT 3.970 195.350 4.330 195.380 ;
        RECT 155.710 195.350 156.070 195.380 ;
        RECT 4.295 195.020 4.655 195.050 ;
        RECT 114.345 195.020 114.725 195.070 ;
        RECT 155.385 195.020 155.745 195.050 ;
        RECT 4.295 194.720 155.750 195.020 ;
        RECT 4.295 194.690 4.655 194.720 ;
        RECT 155.385 194.690 155.745 194.720 ;
        RECT 4.620 194.360 4.980 194.390 ;
        RECT 106.985 194.360 107.365 194.410 ;
        RECT 155.060 194.360 155.420 194.390 ;
        RECT 4.620 194.060 155.425 194.360 ;
        RECT 4.620 194.030 4.980 194.060 ;
        RECT 155.060 194.030 155.420 194.060 ;
        RECT 4.945 193.700 5.305 193.730 ;
        RECT 92.265 193.700 92.645 193.750 ;
        RECT 154.735 193.700 155.095 193.730 ;
        RECT 4.945 193.400 155.100 193.700 ;
        RECT 4.945 193.370 5.305 193.400 ;
        RECT 154.735 193.370 155.095 193.400 ;
        RECT 5.270 193.040 5.630 193.070 ;
        RECT 84.905 193.040 85.285 193.090 ;
        RECT 154.410 193.040 154.770 193.070 ;
        RECT 5.270 192.740 154.775 193.040 ;
        RECT 5.270 192.710 5.630 192.740 ;
        RECT 154.410 192.710 154.770 192.740 ;
        RECT 5.595 192.380 5.955 192.410 ;
        RECT 77.545 192.380 77.925 192.430 ;
        RECT 154.085 192.380 154.445 192.410 ;
        RECT 5.595 192.080 154.450 192.380 ;
        RECT 5.595 192.050 5.955 192.080 ;
        RECT 154.085 192.050 154.445 192.080 ;
        RECT 5.920 191.720 6.280 191.750 ;
        RECT 70.185 191.720 70.565 191.770 ;
        RECT 153.760 191.720 154.120 191.750 ;
        RECT 5.920 191.420 154.125 191.720 ;
        RECT 5.920 191.390 6.280 191.420 ;
        RECT 153.760 191.390 154.120 191.420 ;
        RECT 6.245 191.060 6.605 191.090 ;
        RECT 62.825 191.060 63.205 191.110 ;
        RECT 153.435 191.060 153.795 191.090 ;
        RECT 6.245 190.760 153.800 191.060 ;
        RECT 6.245 190.730 6.605 190.760 ;
        RECT 153.435 190.730 153.795 190.760 ;
        RECT 6.570 190.400 6.930 190.430 ;
        RECT 55.465 190.400 55.845 190.450 ;
        RECT 153.110 190.400 153.470 190.430 ;
        RECT 6.570 190.100 153.475 190.400 ;
        RECT 6.570 190.070 6.930 190.100 ;
        RECT 153.110 190.070 153.470 190.100 ;
        RECT 6.895 189.740 7.255 189.770 ;
        RECT 48.105 189.740 48.485 189.790 ;
        RECT 152.785 189.740 153.145 189.770 ;
        RECT 6.895 189.440 153.150 189.740 ;
        RECT 6.895 189.410 7.255 189.440 ;
        RECT 152.785 189.410 153.145 189.440 ;
        RECT 7.220 189.080 7.580 189.110 ;
        RECT 36.325 189.080 36.705 189.130 ;
        RECT 152.460 189.080 152.820 189.110 ;
        RECT 7.220 188.780 152.825 189.080 ;
        RECT 7.220 188.750 7.580 188.780 ;
        RECT 152.460 188.750 152.820 188.780 ;
        RECT 7.545 188.420 7.905 188.450 ;
        RECT 28.965 188.420 29.345 188.470 ;
        RECT 152.135 188.420 152.495 188.450 ;
        RECT 7.545 188.120 152.500 188.420 ;
        RECT 7.545 188.090 7.905 188.120 ;
        RECT 152.135 188.090 152.495 188.120 ;
        RECT 7.870 187.760 8.230 187.790 ;
        RECT 21.605 187.760 21.985 187.810 ;
        RECT 151.810 187.760 152.170 187.790 ;
        RECT 7.870 187.460 152.175 187.760 ;
        RECT 7.870 187.430 8.230 187.460 ;
        RECT 151.810 187.430 152.170 187.460 ;
        RECT 8.850 161.710 9.850 163.210 ;
        RECT 150.190 159.450 151.190 161.050 ;
        RECT 1.000 157.635 11.240 158.485 ;
        RECT 10.200 157.435 11.240 157.635 ;
        RECT 25.330 157.445 26.360 158.475 ;
        RECT 133.625 157.440 134.655 158.470 ;
        RECT 148.765 157.625 159.040 158.475 ;
        RECT 148.765 157.425 149.840 157.625 ;
        RECT 7.870 156.610 16.085 156.960 ;
        RECT 16.400 156.590 17.055 156.980 ;
        RECT 146.320 156.580 146.975 156.970 ;
        RECT 147.290 156.600 152.190 156.950 ;
        RECT 8.850 151.710 9.850 153.210 ;
        RECT 150.190 149.450 151.190 151.050 ;
        RECT 1.000 147.635 11.240 148.485 ;
        RECT 10.200 147.435 11.240 147.635 ;
        RECT 25.330 147.445 26.360 148.475 ;
        RECT 133.625 147.440 134.655 148.470 ;
        RECT 148.765 147.625 159.040 148.475 ;
        RECT 148.765 147.425 149.840 147.625 ;
        RECT 7.525 146.610 16.085 146.960 ;
        RECT 16.400 146.590 17.055 146.980 ;
        RECT 146.320 146.580 146.975 146.970 ;
        RECT 147.290 146.600 152.515 146.950 ;
        RECT 8.850 141.710 9.850 143.210 ;
        RECT 150.190 139.450 151.190 141.050 ;
        RECT 1.000 137.635 11.240 138.485 ;
        RECT 10.200 137.435 11.240 137.635 ;
        RECT 25.330 137.445 26.360 138.475 ;
        RECT 133.625 137.440 134.655 138.470 ;
        RECT 148.765 137.625 159.040 138.475 ;
        RECT 148.765 137.425 149.840 137.625 ;
        RECT 7.245 136.610 16.085 136.960 ;
        RECT 16.400 136.590 17.055 136.980 ;
        RECT 146.320 136.580 146.975 136.970 ;
        RECT 147.290 136.600 152.840 136.950 ;
        RECT 8.850 131.710 9.850 133.210 ;
        RECT 150.190 129.450 151.190 131.050 ;
        RECT 1.000 127.635 11.240 128.485 ;
        RECT 10.200 127.435 11.240 127.635 ;
        RECT 25.330 127.445 26.360 128.475 ;
        RECT 133.625 127.440 134.655 128.470 ;
        RECT 148.765 127.625 159.040 128.475 ;
        RECT 148.765 127.425 149.840 127.625 ;
        RECT 6.920 126.610 16.085 126.960 ;
        RECT 16.400 126.590 17.055 126.980 ;
        RECT 146.320 126.580 146.975 126.970 ;
        RECT 147.290 126.600 153.165 126.950 ;
        RECT 8.850 121.710 9.850 123.210 ;
        RECT 150.190 119.450 151.190 121.050 ;
        RECT 1.000 117.635 11.240 118.485 ;
        RECT 10.200 117.435 11.240 117.635 ;
        RECT 25.330 117.445 26.360 118.475 ;
        RECT 133.625 117.440 134.655 118.470 ;
        RECT 148.765 117.625 159.040 118.475 ;
        RECT 148.765 117.425 149.840 117.625 ;
        RECT 6.550 116.610 16.085 116.960 ;
        RECT 16.400 116.590 17.055 116.980 ;
        RECT 146.320 116.580 146.975 116.970 ;
        RECT 147.290 116.600 153.490 116.950 ;
        RECT 8.850 111.710 9.850 113.210 ;
        RECT 150.190 109.450 151.190 111.050 ;
        RECT 1.000 107.635 11.240 108.485 ;
        RECT 10.200 107.435 11.240 107.635 ;
        RECT 25.330 107.445 26.360 108.475 ;
        RECT 133.625 107.440 134.655 108.470 ;
        RECT 148.765 107.625 159.040 108.475 ;
        RECT 148.765 107.425 149.840 107.625 ;
        RECT 6.270 106.610 16.085 106.960 ;
        RECT 16.400 106.590 17.055 106.980 ;
        RECT 146.320 106.580 146.975 106.970 ;
        RECT 147.290 106.600 153.815 106.950 ;
        RECT 8.850 101.710 9.850 103.210 ;
        RECT 150.190 99.450 151.190 101.050 ;
        RECT 1.000 97.635 11.240 98.485 ;
        RECT 10.200 97.435 11.240 97.635 ;
        RECT 25.330 97.445 26.360 98.475 ;
        RECT 133.625 97.440 134.655 98.470 ;
        RECT 148.765 97.625 159.040 98.475 ;
        RECT 148.765 97.425 149.840 97.625 ;
        RECT 5.900 96.610 16.085 96.960 ;
        RECT 16.400 96.590 17.055 96.980 ;
        RECT 146.320 96.580 146.975 96.970 ;
        RECT 147.290 96.600 154.140 96.950 ;
        RECT 8.850 91.710 9.850 93.210 ;
        RECT 150.190 89.450 151.190 91.050 ;
        RECT 1.000 87.635 11.240 88.485 ;
        RECT 10.200 87.435 11.240 87.635 ;
        RECT 25.330 87.445 26.360 88.475 ;
        RECT 133.625 87.440 134.655 88.470 ;
        RECT 148.765 87.625 159.040 88.475 ;
        RECT 148.765 87.425 149.840 87.625 ;
        RECT 5.575 86.610 16.085 86.960 ;
        RECT 16.400 86.590 17.055 86.980 ;
        RECT 146.320 86.580 146.975 86.970 ;
        RECT 147.290 86.600 154.465 86.950 ;
        RECT 8.850 81.710 9.850 83.210 ;
        RECT 150.190 79.450 151.190 81.050 ;
        RECT 1.000 77.635 11.240 78.485 ;
        RECT 10.200 77.435 11.240 77.635 ;
        RECT 25.330 77.445 26.360 78.475 ;
        RECT 133.625 77.440 134.655 78.470 ;
        RECT 148.765 77.625 159.040 78.475 ;
        RECT 148.765 77.425 149.840 77.625 ;
        RECT 5.250 76.610 16.085 76.960 ;
        RECT 16.400 76.590 17.055 76.980 ;
        RECT 146.320 76.580 146.975 76.970 ;
        RECT 147.290 76.600 154.790 76.950 ;
        RECT 8.850 71.710 9.850 73.210 ;
        RECT 150.190 69.450 151.190 71.050 ;
        RECT 1.000 67.635 11.240 68.485 ;
        RECT 10.200 67.435 11.240 67.635 ;
        RECT 25.330 67.445 26.360 68.475 ;
        RECT 133.625 67.440 134.655 68.470 ;
        RECT 148.765 67.625 159.040 68.475 ;
        RECT 148.765 67.425 149.840 67.625 ;
        RECT 4.925 66.610 16.085 66.960 ;
        RECT 16.400 66.590 17.055 66.980 ;
        RECT 146.320 66.580 146.975 66.970 ;
        RECT 147.290 66.600 155.115 66.950 ;
        RECT 8.850 61.710 9.850 63.210 ;
        RECT 150.190 59.450 151.190 61.050 ;
        RECT 1.000 57.635 11.240 58.485 ;
        RECT 10.200 57.435 11.240 57.635 ;
        RECT 25.330 57.445 26.360 58.475 ;
        RECT 133.625 57.440 134.655 58.470 ;
        RECT 148.765 57.625 159.040 58.475 ;
        RECT 148.765 57.425 149.840 57.625 ;
        RECT 4.600 56.610 16.085 56.960 ;
        RECT 16.400 56.590 17.055 56.980 ;
        RECT 146.320 56.580 146.975 56.970 ;
        RECT 147.290 56.600 155.440 56.950 ;
        RECT 8.850 51.710 9.850 53.210 ;
        RECT 150.190 49.450 151.190 51.050 ;
        RECT 1.000 47.635 11.240 48.485 ;
        RECT 10.200 47.435 11.240 47.635 ;
        RECT 25.330 47.445 26.360 48.475 ;
        RECT 133.625 47.440 134.655 48.470 ;
        RECT 148.765 47.625 159.040 48.475 ;
        RECT 148.765 47.425 149.840 47.625 ;
        RECT 4.275 46.610 16.085 46.960 ;
        RECT 16.400 46.590 17.055 46.980 ;
        RECT 146.320 46.580 146.975 46.970 ;
        RECT 147.290 46.600 155.765 46.950 ;
        RECT 8.850 41.710 9.850 43.210 ;
        RECT 150.190 39.450 151.190 41.050 ;
        RECT 1.000 37.635 11.240 38.485 ;
        RECT 10.200 37.435 11.240 37.635 ;
        RECT 25.330 37.445 26.360 38.475 ;
        RECT 133.625 37.440 134.655 38.470 ;
        RECT 148.765 37.625 159.040 38.475 ;
        RECT 148.765 37.425 149.840 37.625 ;
        RECT 3.940 36.610 16.085 36.960 ;
        RECT 16.400 36.590 17.055 36.980 ;
        RECT 146.320 36.580 146.975 36.970 ;
        RECT 147.290 36.600 156.090 36.950 ;
        RECT 8.850 31.710 9.850 33.210 ;
        RECT 150.190 29.450 151.190 31.050 ;
        RECT 1.000 27.635 11.240 28.485 ;
        RECT 10.200 27.435 11.240 27.635 ;
        RECT 25.330 27.445 26.360 28.475 ;
        RECT 133.625 27.440 134.655 28.470 ;
        RECT 148.765 27.625 159.040 28.475 ;
        RECT 148.765 27.425 149.840 27.625 ;
        RECT 3.625 26.610 16.085 26.960 ;
        RECT 16.400 26.590 17.055 26.980 ;
        RECT 146.320 26.580 146.975 26.970 ;
        RECT 147.290 26.600 156.415 26.950 ;
        RECT 8.850 21.710 9.850 23.210 ;
        RECT 150.190 19.450 151.190 21.050 ;
        RECT 1.000 17.635 11.240 18.485 ;
        RECT 10.200 17.435 11.240 17.635 ;
        RECT 25.330 17.445 26.360 18.475 ;
        RECT 133.625 17.440 134.655 18.470 ;
        RECT 148.765 17.625 159.040 18.475 ;
        RECT 148.765 17.425 149.840 17.625 ;
        RECT 3.290 16.610 16.085 16.960 ;
        RECT 16.400 16.590 17.055 16.980 ;
        RECT 146.320 16.580 146.975 16.970 ;
        RECT 147.290 16.600 156.740 16.950 ;
        RECT 8.850 11.710 9.850 13.210 ;
        RECT 150.190 9.450 151.190 11.050 ;
        RECT 1.000 7.635 11.240 8.485 ;
        RECT 10.200 7.435 11.240 7.635 ;
        RECT 25.330 7.445 26.360 8.475 ;
        RECT 133.625 7.440 134.655 8.470 ;
        RECT 148.765 7.625 159.040 8.475 ;
        RECT 148.765 7.425 149.840 7.625 ;
        RECT 2.975 6.610 16.085 6.960 ;
        RECT 16.400 6.590 17.055 6.980 ;
        RECT 146.320 6.580 146.975 6.970 ;
        RECT 147.290 6.600 157.065 6.950 ;
        RECT 134.280 5.150 151.190 5.200 ;
        RECT 134.280 4.250 151.200 5.150 ;
        RECT 134.280 4.200 151.190 4.250 ;
        RECT 123.450 2.200 124.450 3.200 ;
        RECT 123.450 1.200 157.360 2.200 ;
      LAYER met4 ;
        RECT 3.990 222.775 4.290 224.760 ;
        RECT 7.670 222.775 7.970 224.760 ;
        RECT 11.350 222.775 11.650 224.760 ;
        RECT 15.030 222.775 15.330 224.760 ;
        RECT 18.710 222.775 19.010 224.760 ;
        RECT 22.390 224.135 22.690 224.760 ;
        RECT 22.375 223.805 22.705 224.135 ;
        RECT 3.975 222.445 4.305 222.775 ;
        RECT 7.655 222.445 7.985 222.775 ;
        RECT 11.335 222.445 11.665 222.775 ;
        RECT 15.015 222.445 15.345 222.775 ;
        RECT 18.695 222.445 19.025 222.775 ;
        RECT 6.735 205.445 7.065 205.775 ;
        RECT 14.095 205.445 14.425 205.775 ;
        RECT 6.750 200.320 7.050 205.445 ;
        RECT 14.110 200.320 14.410 205.445 ;
        RECT 21.395 201.040 22.995 223.280 ;
        RECT 26.070 222.775 26.370 224.760 ;
        RECT 29.750 222.775 30.050 224.760 ;
        RECT 26.055 222.445 26.385 222.775 ;
        RECT 29.735 222.445 30.065 222.775 ;
        RECT 33.430 208.495 33.730 224.760 ;
        RECT 37.110 211.215 37.410 224.760 ;
        RECT 40.790 224.120 41.090 224.760 ;
        RECT 39.870 223.820 41.090 224.120 ;
        RECT 37.095 210.885 37.425 211.215 ;
        RECT 39.870 210.535 40.170 223.820 ;
        RECT 39.855 210.205 40.185 210.535 ;
        RECT 44.470 209.175 44.770 224.760 ;
        RECT 48.150 223.455 48.450 224.760 ;
        RECT 48.135 223.125 48.465 223.455 ;
        RECT 51.830 209.855 52.130 224.760 ;
        RECT 51.815 209.525 52.145 209.855 ;
        RECT 44.455 208.845 44.785 209.175 ;
        RECT 33.415 208.165 33.745 208.495 ;
        RECT 23.295 207.485 23.625 207.815 ;
        RECT 23.310 200.320 23.610 207.485 ;
        RECT 55.510 207.135 55.810 224.760 ;
        RECT 55.495 206.805 55.825 207.135 ;
        RECT 59.190 206.455 59.490 224.760 ;
        RECT 48.135 206.125 48.465 206.455 ;
        RECT 59.175 206.125 59.505 206.455 ;
        RECT 28.815 205.445 29.145 205.775 ;
        RECT 36.175 205.445 36.505 205.775 ;
        RECT 6.750 200.020 7.225 200.320 ;
        RECT 14.110 200.020 14.585 200.320 ;
        RECT 6.925 199.020 7.225 200.020 ;
        RECT 14.285 199.020 14.585 200.020 ;
        RECT 21.645 200.020 23.610 200.320 ;
        RECT 28.830 200.320 29.130 205.445 ;
        RECT 36.190 200.320 36.490 205.445 ;
        RECT 28.830 200.020 29.305 200.320 ;
        RECT 36.190 200.020 36.665 200.320 ;
        RECT 21.645 199.020 21.945 200.020 ;
        RECT 29.005 199.020 29.305 200.020 ;
        RECT 36.365 199.020 36.665 200.020 ;
        RECT 48.150 199.020 48.450 206.125 ;
        RECT 55.495 205.445 55.825 205.775 ;
        RECT 55.510 199.020 55.810 205.445 ;
        RECT 60.265 201.040 61.865 223.280 ;
        RECT 62.870 222.775 63.170 224.760 ;
        RECT 62.855 222.445 63.185 222.775 ;
        RECT 66.550 211.895 66.850 224.760 ;
        RECT 70.230 219.375 70.530 224.760 ;
        RECT 70.215 219.045 70.545 219.375 ;
        RECT 73.910 216.655 74.210 224.760 ;
        RECT 77.590 222.095 77.890 224.760 ;
        RECT 81.270 224.135 81.570 224.760 ;
        RECT 81.255 223.805 81.585 224.135 ;
        RECT 77.575 221.765 77.905 222.095 ;
        RECT 73.895 216.325 74.225 216.655 ;
        RECT 66.535 211.565 66.865 211.895 ;
        RECT 77.575 205.445 77.905 205.775 ;
        RECT 70.215 200.685 70.545 201.015 ;
        RECT 62.855 200.005 63.185 200.335 ;
        RECT 62.870 199.020 63.170 200.005 ;
        RECT 70.230 199.020 70.530 200.685 ;
        RECT 77.590 199.020 77.890 205.445 ;
        RECT 79.700 201.040 81.300 223.280 ;
        RECT 84.950 222.095 85.250 224.760 ;
        RECT 88.630 224.135 88.930 224.760 ;
        RECT 121.750 224.135 122.050 224.760 ;
        RECT 88.615 223.805 88.945 224.135 ;
        RECT 121.735 223.805 122.065 224.135 ;
        RECT 125.430 223.455 125.730 224.760 ;
        RECT 132.790 223.455 133.090 224.760 ;
        RECT 136.470 223.455 136.770 224.760 ;
        RECT 84.935 221.765 85.265 222.095 ;
        RECT 92.295 205.445 92.625 205.775 ;
        RECT 107.015 205.445 107.345 205.775 ;
        RECT 114.375 205.445 114.705 205.775 ;
        RECT 84.935 200.005 85.265 200.335 ;
        RECT 84.950 199.020 85.250 200.005 ;
        RECT 92.310 199.020 92.610 205.445 ;
        RECT 107.030 199.020 107.330 205.445 ;
        RECT 114.390 199.020 114.690 205.445 ;
        RECT 118.570 201.040 120.170 223.280 ;
        RECT 125.415 223.125 125.745 223.455 ;
        RECT 132.775 223.125 133.105 223.455 ;
        RECT 136.455 223.125 136.785 223.455 ;
        RECT 121.735 205.445 122.065 205.775 ;
        RECT 129.095 205.445 129.425 205.775 ;
        RECT 121.750 199.020 122.050 205.445 ;
        RECT 129.110 199.020 129.410 205.445 ;
        RECT 136.455 201.365 136.785 201.695 ;
        RECT 136.470 199.020 136.770 201.365 ;
        RECT 138.005 201.040 139.605 223.280 ;
        RECT 140.150 220.735 140.450 224.760 ;
        RECT 140.135 220.405 140.465 220.735 ;
        RECT 143.830 219.375 144.130 224.760 ;
        RECT 147.510 220.735 147.810 224.760 ;
        RECT 147.495 220.405 147.825 220.735 ;
        RECT 143.815 219.045 144.145 219.375 ;
        RECT 151.190 211.215 151.490 224.760 ;
        RECT 154.870 220.055 155.170 224.760 ;
        RECT 158.550 224.120 158.850 224.760 ;
        RECT 156.710 223.820 158.850 224.120 ;
        RECT 154.855 219.725 155.185 220.055 ;
        RECT 151.175 210.885 151.505 211.215 ;
        RECT 156.710 209.175 157.010 223.820 ;
        RECT 156.695 208.845 157.025 209.175 ;
        RECT 151.175 205.445 151.505 205.775 ;
        RECT 143.815 200.685 144.145 201.015 ;
        RECT 143.830 199.020 144.130 200.685 ;
        RECT 151.190 199.020 151.490 205.445 ;
        RECT 6.880 198.625 6.925 199.015 ;
        RECT 7.225 198.625 7.270 199.015 ;
        RECT 14.240 198.625 14.285 199.015 ;
        RECT 14.585 198.625 14.630 199.015 ;
        RECT 151.145 198.020 151.190 198.370 ;
        RECT 151.490 198.020 151.525 198.370 ;
        RECT 21.645 187.810 21.945 198.020 ;
        RECT 29.005 188.470 29.305 198.020 ;
        RECT 36.365 189.130 36.665 198.020 ;
        RECT 48.150 189.790 48.450 198.020 ;
        RECT 55.510 190.450 55.810 198.020 ;
        RECT 62.870 191.110 63.170 198.020 ;
        RECT 70.230 191.770 70.530 198.020 ;
        RECT 77.590 192.430 77.890 198.020 ;
        RECT 84.950 193.090 85.250 198.020 ;
        RECT 92.310 193.750 92.610 198.020 ;
        RECT 107.030 194.410 107.330 198.020 ;
        RECT 114.390 195.070 114.690 198.020 ;
        RECT 121.750 195.730 122.050 198.020 ;
        RECT 129.110 196.390 129.410 198.020 ;
        RECT 136.470 197.050 136.770 198.020 ;
        RECT 143.830 197.710 144.130 198.020 ;
        RECT 143.785 197.360 144.165 197.710 ;
        RECT 136.425 196.700 136.805 197.050 ;
        RECT 129.065 196.040 129.445 196.390 ;
        RECT 121.705 195.380 122.085 195.730 ;
        RECT 114.345 194.720 114.725 195.070 ;
        RECT 106.985 194.060 107.365 194.410 ;
        RECT 92.265 193.400 92.645 193.750 ;
        RECT 84.905 192.740 85.285 193.090 ;
        RECT 77.545 192.080 77.925 192.430 ;
        RECT 70.185 191.420 70.565 191.770 ;
        RECT 62.825 190.760 63.205 191.110 ;
        RECT 55.465 190.100 55.845 190.450 ;
        RECT 48.105 189.440 48.485 189.790 ;
        RECT 36.325 188.780 36.705 189.130 ;
        RECT 28.965 188.120 29.345 188.470 ;
        RECT 21.605 187.460 21.985 187.810 ;
        RECT 8.200 158.485 8.500 166.500 ;
        RECT 2.600 157.635 8.500 158.485 ;
        RECT 8.200 148.485 8.500 157.635 ;
        RECT 2.600 147.635 8.500 148.485 ;
        RECT 8.200 138.485 8.500 147.635 ;
        RECT 2.600 137.635 8.500 138.485 ;
        RECT 8.200 128.485 8.500 137.635 ;
        RECT 2.600 127.635 8.500 128.485 ;
        RECT 8.200 118.485 8.500 127.635 ;
        RECT 2.600 117.635 8.500 118.485 ;
        RECT 8.200 108.485 8.500 117.635 ;
        RECT 2.600 107.635 8.500 108.485 ;
        RECT 8.200 98.485 8.500 107.635 ;
        RECT 2.600 97.635 8.500 98.485 ;
        RECT 8.200 88.485 8.500 97.635 ;
        RECT 2.600 87.635 8.500 88.485 ;
        RECT 8.200 78.485 8.500 87.635 ;
        RECT 2.600 77.635 8.500 78.485 ;
        RECT 8.200 68.485 8.500 77.635 ;
        RECT 2.600 67.635 8.500 68.485 ;
        RECT 8.200 58.485 8.500 67.635 ;
        RECT 2.600 57.635 8.500 58.485 ;
        RECT 8.200 48.485 8.500 57.635 ;
        RECT 2.600 47.635 8.500 48.485 ;
        RECT 8.200 38.485 8.500 47.635 ;
        RECT 2.600 37.635 8.500 38.485 ;
        RECT 8.200 28.485 8.500 37.635 ;
        RECT 2.600 27.635 8.500 28.485 ;
        RECT 8.200 18.485 8.500 27.635 ;
        RECT 2.600 17.635 8.500 18.485 ;
        RECT 8.200 8.485 8.500 17.635 ;
        RECT 2.600 7.635 8.500 8.485 ;
        RECT 8.200 6.000 8.500 7.635 ;
        RECT 8.850 3.200 9.850 166.500 ;
        RECT 10.200 158.460 10.500 166.500 ;
        RECT 149.540 158.475 149.840 166.490 ;
        RECT 10.195 157.460 10.550 158.460 ;
        RECT 25.345 157.460 40.830 158.460 ;
        RECT 10.200 148.460 10.500 157.460 ;
        RECT 15.635 156.610 17.040 156.960 ;
        RECT 26.440 148.460 27.090 157.460 ;
        RECT 100.735 157.455 134.640 158.455 ;
        RECT 10.195 147.460 10.550 148.460 ;
        RECT 25.345 147.460 27.090 148.460 ;
        RECT 10.200 138.460 10.500 147.460 ;
        RECT 15.635 146.610 17.040 146.960 ;
        RECT 26.440 138.460 27.090 147.460 ;
        RECT 10.195 137.460 10.550 138.460 ;
        RECT 25.345 137.460 27.090 138.460 ;
        RECT 10.200 128.460 10.500 137.460 ;
        RECT 15.635 136.610 17.040 136.960 ;
        RECT 26.440 128.460 27.090 137.460 ;
        RECT 10.195 127.460 10.550 128.460 ;
        RECT 25.345 127.460 27.090 128.460 ;
        RECT 10.200 118.460 10.500 127.460 ;
        RECT 15.635 126.610 17.040 126.960 ;
        RECT 26.440 118.460 27.090 127.460 ;
        RECT 10.195 117.460 10.550 118.460 ;
        RECT 25.345 117.460 27.090 118.460 ;
        RECT 10.200 108.460 10.500 117.460 ;
        RECT 15.635 116.610 17.040 116.960 ;
        RECT 26.440 108.460 27.090 117.460 ;
        RECT 10.195 107.460 10.550 108.460 ;
        RECT 25.345 107.460 27.090 108.460 ;
        RECT 10.200 98.460 10.500 107.460 ;
        RECT 15.635 106.610 17.040 106.960 ;
        RECT 26.440 98.460 27.090 107.460 ;
        RECT 10.195 97.460 10.550 98.460 ;
        RECT 25.345 97.460 27.090 98.460 ;
        RECT 10.200 88.460 10.500 97.460 ;
        RECT 15.635 96.610 17.040 96.960 ;
        RECT 26.440 88.460 27.090 97.460 ;
        RECT 10.195 87.460 10.550 88.460 ;
        RECT 25.345 87.460 27.090 88.460 ;
        RECT 10.200 78.460 10.500 87.460 ;
        RECT 15.635 86.610 17.040 86.960 ;
        RECT 26.440 78.460 27.090 87.460 ;
        RECT 10.195 77.460 10.550 78.460 ;
        RECT 25.345 77.460 27.090 78.460 ;
        RECT 10.200 68.460 10.500 77.460 ;
        RECT 15.635 76.610 17.040 76.960 ;
        RECT 26.440 68.460 27.090 77.460 ;
        RECT 10.195 67.460 10.550 68.460 ;
        RECT 25.345 67.460 27.090 68.460 ;
        RECT 10.200 58.460 10.500 67.460 ;
        RECT 15.635 66.610 17.040 66.960 ;
        RECT 26.440 58.460 27.090 67.460 ;
        RECT 10.195 57.460 10.550 58.460 ;
        RECT 25.345 57.460 27.090 58.460 ;
        RECT 10.200 48.460 10.500 57.460 ;
        RECT 15.635 56.610 17.040 56.960 ;
        RECT 26.440 48.460 27.090 57.460 ;
        RECT 10.195 47.460 10.550 48.460 ;
        RECT 25.345 47.460 27.090 48.460 ;
        RECT 10.200 38.460 10.500 47.460 ;
        RECT 15.635 46.610 17.040 46.960 ;
        RECT 26.440 38.460 27.090 47.460 ;
        RECT 10.195 37.460 10.550 38.460 ;
        RECT 25.345 37.460 27.090 38.460 ;
        RECT 10.200 28.460 10.500 37.460 ;
        RECT 15.635 36.610 17.040 36.960 ;
        RECT 26.440 28.460 27.090 37.460 ;
        RECT 10.195 27.460 10.550 28.460 ;
        RECT 25.345 27.460 27.090 28.460 ;
        RECT 10.200 18.460 10.500 27.460 ;
        RECT 15.635 26.610 17.040 26.960 ;
        RECT 26.440 18.460 27.090 27.460 ;
        RECT 10.195 17.460 10.550 18.460 ;
        RECT 25.345 17.460 27.090 18.460 ;
        RECT 10.200 8.460 10.500 17.460 ;
        RECT 15.635 16.610 17.040 16.960 ;
        RECT 26.440 8.460 27.090 17.460 ;
        RECT 132.890 148.455 133.540 157.455 ;
        RECT 148.765 157.425 149.840 158.475 ;
        RECT 146.320 156.600 147.750 156.950 ;
        RECT 149.540 148.475 149.840 157.425 ;
        RECT 132.890 147.455 134.640 148.455 ;
        RECT 132.890 138.455 133.540 147.455 ;
        RECT 148.765 147.425 149.840 148.475 ;
        RECT 146.320 146.600 147.750 146.950 ;
        RECT 149.540 138.475 149.840 147.425 ;
        RECT 132.890 137.455 134.640 138.455 ;
        RECT 132.890 128.455 133.540 137.455 ;
        RECT 148.765 137.425 149.840 138.475 ;
        RECT 146.320 136.600 147.750 136.950 ;
        RECT 149.540 128.475 149.840 137.425 ;
        RECT 132.890 127.455 134.640 128.455 ;
        RECT 132.890 118.455 133.540 127.455 ;
        RECT 148.765 127.425 149.840 128.475 ;
        RECT 146.320 126.600 147.750 126.950 ;
        RECT 149.540 118.475 149.840 127.425 ;
        RECT 132.890 117.455 134.640 118.455 ;
        RECT 132.890 108.455 133.540 117.455 ;
        RECT 148.765 117.425 149.840 118.475 ;
        RECT 146.320 116.600 147.750 116.950 ;
        RECT 149.540 108.475 149.840 117.425 ;
        RECT 132.890 107.455 134.640 108.455 ;
        RECT 132.890 98.455 133.540 107.455 ;
        RECT 148.765 107.425 149.840 108.475 ;
        RECT 146.320 106.600 147.750 106.950 ;
        RECT 149.540 98.475 149.840 107.425 ;
        RECT 132.890 97.455 134.640 98.455 ;
        RECT 132.890 88.455 133.540 97.455 ;
        RECT 148.765 97.425 149.840 98.475 ;
        RECT 146.320 96.600 147.750 96.950 ;
        RECT 149.540 88.475 149.840 97.425 ;
        RECT 132.890 87.455 134.640 88.455 ;
        RECT 132.890 78.455 133.540 87.455 ;
        RECT 148.765 87.425 149.840 88.475 ;
        RECT 146.320 86.600 147.750 86.950 ;
        RECT 149.540 78.475 149.840 87.425 ;
        RECT 132.890 77.455 134.640 78.455 ;
        RECT 132.890 68.455 133.540 77.455 ;
        RECT 148.765 77.425 149.840 78.475 ;
        RECT 146.320 76.600 147.750 76.950 ;
        RECT 149.540 68.475 149.840 77.425 ;
        RECT 132.890 67.455 134.640 68.455 ;
        RECT 132.890 58.455 133.540 67.455 ;
        RECT 148.765 67.425 149.840 68.475 ;
        RECT 146.320 66.600 147.750 66.950 ;
        RECT 149.540 58.475 149.840 67.425 ;
        RECT 132.890 57.455 134.640 58.455 ;
        RECT 132.890 48.455 133.540 57.455 ;
        RECT 148.765 57.425 149.840 58.475 ;
        RECT 146.320 56.600 147.750 56.950 ;
        RECT 149.540 48.475 149.840 57.425 ;
        RECT 132.890 47.455 134.640 48.455 ;
        RECT 132.890 38.455 133.540 47.455 ;
        RECT 148.765 47.425 149.840 48.475 ;
        RECT 146.320 46.600 147.750 46.950 ;
        RECT 149.540 38.475 149.840 47.425 ;
        RECT 132.890 37.455 134.640 38.455 ;
        RECT 132.890 28.455 133.540 37.455 ;
        RECT 148.765 37.425 149.840 38.475 ;
        RECT 146.320 36.600 147.750 36.950 ;
        RECT 149.540 28.475 149.840 37.425 ;
        RECT 132.890 27.455 134.640 28.455 ;
        RECT 132.890 18.455 133.540 27.455 ;
        RECT 148.765 27.425 149.840 28.475 ;
        RECT 146.320 26.600 147.750 26.950 ;
        RECT 149.540 18.475 149.840 27.425 ;
        RECT 132.890 17.455 134.640 18.455 ;
        RECT 10.195 7.460 10.550 8.460 ;
        RECT 25.345 7.460 40.830 8.460 ;
        RECT 132.890 8.455 133.540 17.455 ;
        RECT 148.765 17.425 149.840 18.475 ;
        RECT 146.320 16.600 147.750 16.950 ;
        RECT 149.540 8.475 149.840 17.425 ;
        RECT 10.200 6.000 10.500 7.460 ;
        RECT 26.440 7.455 27.090 7.460 ;
        RECT 100.735 7.455 134.640 8.455 ;
        RECT 148.765 7.425 149.840 8.475 ;
        RECT 15.635 6.610 17.040 6.960 ;
        RECT 146.320 6.600 147.750 6.950 ;
        RECT 149.540 5.990 149.840 7.425 ;
        RECT 8.850 2.200 124.450 3.200 ;
        RECT 134.280 1.000 135.280 5.200 ;
        RECT 150.190 4.200 151.190 166.490 ;
        RECT 151.540 158.475 151.840 166.490 ;
        RECT 151.540 157.625 157.440 158.475 ;
        RECT 151.540 148.475 151.840 157.625 ;
        RECT 151.540 147.625 157.440 148.475 ;
        RECT 151.540 138.475 151.840 147.625 ;
        RECT 151.540 137.625 157.440 138.475 ;
        RECT 151.540 128.475 151.840 137.625 ;
        RECT 151.540 127.625 157.440 128.475 ;
        RECT 151.540 118.475 151.840 127.625 ;
        RECT 151.540 117.625 157.440 118.475 ;
        RECT 151.540 108.475 151.840 117.625 ;
        RECT 151.540 107.625 157.440 108.475 ;
        RECT 151.540 98.475 151.840 107.625 ;
        RECT 151.540 97.625 157.440 98.475 ;
        RECT 151.540 88.475 151.840 97.625 ;
        RECT 151.540 87.625 157.440 88.475 ;
        RECT 151.540 78.475 151.840 87.625 ;
        RECT 151.540 77.625 157.440 78.475 ;
        RECT 151.540 68.475 151.840 77.625 ;
        RECT 151.540 67.625 157.440 68.475 ;
        RECT 151.540 58.475 151.840 67.625 ;
        RECT 151.540 57.625 157.440 58.475 ;
        RECT 151.540 48.475 151.840 57.625 ;
        RECT 151.540 47.625 157.440 48.475 ;
        RECT 151.540 38.475 151.840 47.625 ;
        RECT 151.540 37.625 157.440 38.475 ;
        RECT 151.540 28.475 151.840 37.625 ;
        RECT 151.540 27.625 157.440 28.475 ;
        RECT 151.540 18.475 151.840 27.625 ;
        RECT 151.540 17.625 157.440 18.475 ;
        RECT 151.540 8.475 151.840 17.625 ;
        RECT 151.540 7.625 157.440 8.475 ;
        RECT 151.540 5.990 151.840 7.625 ;
        RECT 134.280 0.000 134.330 1.000 ;
        RECT 135.230 0.000 135.280 1.000 ;
        RECT 156.360 1.000 157.360 2.200 ;
        RECT 156.360 0.000 156.410 1.000 ;
        RECT 157.310 0.000 157.360 1.000 ;
  END
END tt_um_dlmiles_schmitt_playground
END LIBRARY

