magic
tech sky130A
magscale 1 2
timestamp 1717265471
<< locali >>
rect 1407 2033 3770 2100
rect 1407 2015 1990 2033
rect 1407 489 1863 2015
rect 1907 532 1990 2015
rect 2120 532 3310 533
rect 1907 492 3310 532
rect 1407 294 1423 489
rect 3247 294 3310 492
rect 1407 68 3310 294
rect 3595 68 3770 2033
rect 1407 0 3770 68
rect 3805 1975 5070 2100
rect 3805 1612 4983 1975
rect 3805 73 3980 1612
rect 4818 539 4983 1612
rect 4265 518 4490 533
rect 4265 349 4351 518
rect 4423 349 4490 518
rect 4265 73 4490 349
rect 3805 52 4490 73
rect 4818 294 4833 539
rect 5027 489 5070 1975
rect 5054 294 5070 489
rect 4818 52 4983 294
rect 3805 19 4983 52
rect 5027 19 5070 294
rect 3805 0 5070 19
<< viali >>
rect 1863 492 1907 2015
rect 1863 489 3247 492
rect 1423 294 3247 489
rect 4983 539 5027 1975
rect 4351 349 4423 518
rect 4833 489 5027 539
rect 4833 294 5054 489
rect 4983 19 5027 294
<< metal1 >>
rect 1850 2015 1920 2097
rect 1850 499 1863 2015
rect 1410 492 1863 499
rect 1907 499 1920 2015
rect 2120 1917 3740 1977
rect 2064 1432 2110 1876
rect 2055 1152 2065 1432
rect 2137 1152 2147 1432
rect 2064 686 2110 1152
rect 2192 992 2238 1876
rect 2320 1432 2366 1876
rect 2310 1152 2320 1432
rect 2392 1152 2402 1432
rect 2185 712 2195 992
rect 2267 712 2277 992
rect 2192 686 2238 712
rect 2320 686 2366 1152
rect 2448 992 2494 1876
rect 2576 1432 2622 1876
rect 2565 1152 2575 1432
rect 2647 1152 2657 1432
rect 2443 712 2453 992
rect 2525 712 2535 992
rect 2448 686 2494 712
rect 2576 686 2622 1152
rect 2704 992 2750 1876
rect 2832 1432 2878 1876
rect 2820 1152 2830 1432
rect 2902 1152 2912 1432
rect 2698 712 2708 992
rect 2780 712 2790 992
rect 2704 686 2750 712
rect 2832 686 2878 1152
rect 2960 992 3006 1876
rect 3088 1432 3134 1876
rect 3075 1152 3085 1432
rect 3157 1152 3167 1432
rect 2953 712 2963 992
rect 3035 712 3045 992
rect 2960 686 3006 712
rect 3088 686 3134 1152
rect 3216 992 3262 1876
rect 3344 1432 3390 1876
rect 3330 1152 3340 1432
rect 3412 1152 3422 1432
rect 3208 712 3218 992
rect 3290 712 3300 992
rect 3216 686 3262 712
rect 3344 686 3390 1152
rect 3472 992 3518 1876
rect 3660 1682 3740 1917
rect 4970 1975 5040 2096
rect 4870 1684 4940 1692
rect 4870 1682 4878 1684
rect 3660 1622 4878 1682
rect 3463 712 3473 992
rect 3545 712 3555 992
rect 3472 686 3518 712
rect 3660 642 3740 1622
rect 4870 1620 4878 1622
rect 4932 1620 4940 1684
rect 4870 1612 4940 1620
rect 4110 1502 4940 1562
rect 4056 1432 4102 1466
rect 4045 1152 4055 1432
rect 4127 1152 4137 1432
rect 4056 678 4102 1152
rect 4184 992 4230 1466
rect 4312 1432 4358 1466
rect 4300 1152 4310 1432
rect 4382 1152 4392 1432
rect 4178 712 4188 992
rect 4260 712 4270 992
rect 4184 678 4230 712
rect 4312 678 4358 1152
rect 4440 992 4486 1466
rect 4568 1432 4614 1466
rect 4555 1152 4565 1432
rect 4637 1152 4647 1432
rect 4433 712 4443 992
rect 4515 712 4525 992
rect 4440 678 4486 712
rect 4568 678 4614 1152
rect 4696 992 4742 1466
rect 4886 1352 4940 1502
rect 4870 1344 4940 1352
rect 4870 1280 4878 1344
rect 4932 1280 4940 1344
rect 4870 1272 4940 1280
rect 4690 712 4700 992
rect 4752 712 4762 992
rect 4696 678 4742 712
rect 4886 642 4940 1272
rect 2120 582 3740 642
rect 1907 492 3260 499
rect 1410 489 1848 492
rect 1410 294 1423 489
rect 3247 294 3260 492
rect 3384 402 3430 414
rect 3472 402 3518 414
rect 3660 402 3740 582
rect 3832 582 4940 642
rect 3363 332 3373 402
rect 3425 332 3435 402
rect 3468 332 3478 402
rect 3530 332 3540 402
rect 3650 332 3660 402
rect 3740 332 3750 402
rect 1410 292 1848 294
rect 1900 292 3260 294
rect 1410 286 3260 292
rect 3384 226 3430 332
rect 3472 226 3518 332
rect 3660 322 3740 332
rect 3120 184 3210 192
rect 3120 130 3128 184
rect 3202 182 3210 184
rect 3832 182 3912 582
rect 4970 552 4983 1975
rect 4334 539 4983 552
rect 4334 518 4833 539
rect 4056 402 4102 406
rect 4144 402 4190 406
rect 4334 404 4351 518
rect 4423 512 4833 518
rect 4423 404 4440 512
rect 4033 332 4043 402
rect 4095 332 4105 402
rect 4138 332 4148 402
rect 4200 332 4210 402
rect 4334 340 4342 404
rect 4432 340 4440 404
rect 4584 402 4630 406
rect 4334 332 4440 340
rect 4555 394 4630 402
rect 4555 340 4563 394
rect 4617 340 4630 394
rect 4555 332 4630 340
rect 4056 218 4102 332
rect 4144 218 4190 332
rect 4584 218 4630 332
rect 4672 402 4718 406
rect 4672 394 4748 402
rect 4672 340 4686 394
rect 4740 340 4748 394
rect 4672 332 4748 340
rect 4672 218 4718 332
rect 4820 294 4833 512
rect 5027 499 5040 1975
rect 5027 492 5067 499
rect 5062 294 5067 492
rect 4820 286 4983 294
rect 3202 132 4147 182
rect 4605 179 4695 183
rect 3202 130 3210 132
rect 3120 122 3210 130
rect 4605 120 4615 179
rect 4685 120 4695 179
rect 4605 119 4695 120
rect 4970 19 4983 286
rect 5027 286 5067 294
rect 5027 19 5040 286
rect 4970 8 5040 19
<< via1 >>
rect 2065 1152 2137 1432
rect 2320 1152 2392 1432
rect 2195 712 2267 992
rect 2575 1152 2647 1432
rect 2453 712 2525 992
rect 2830 1152 2902 1432
rect 2708 712 2780 992
rect 3085 1152 3157 1432
rect 2963 712 3035 992
rect 3340 1152 3412 1432
rect 3218 712 3290 992
rect 3473 712 3545 992
rect 4878 1620 4932 1684
rect 4055 1152 4127 1432
rect 4310 1152 4382 1432
rect 4188 712 4260 992
rect 4565 1152 4637 1432
rect 4443 712 4515 992
rect 4878 1280 4932 1344
rect 4700 712 4752 992
rect 1848 489 1863 492
rect 1863 491 1900 492
rect 1863 489 2041 491
rect 1440 335 1505 489
rect 1848 294 2041 489
rect 3163 342 3247 482
rect 3373 332 3425 402
rect 3478 332 3530 402
rect 3660 332 3740 402
rect 1848 292 1900 294
rect 3128 130 3202 184
rect 4043 332 4095 402
rect 4148 332 4200 402
rect 4342 349 4351 404
rect 4351 349 4423 404
rect 4423 349 4432 404
rect 4342 340 4432 349
rect 4563 340 4617 394
rect 4686 340 4740 394
rect 4878 489 5027 492
rect 5027 489 5062 492
rect 4878 294 5054 489
rect 5054 294 5062 489
rect 4615 120 4685 179
<< metal2 >>
rect 334 0 367 2100
rect 399 0 432 2100
rect 464 0 497 2100
rect 529 0 562 2100
rect 594 0 627 2100
rect 659 0 692 2100
rect 724 0 757 2100
rect 789 0 822 2100
rect 854 0 887 2100
rect 919 0 952 2100
rect 984 0 1017 2100
rect 1049 0 1082 2100
rect 1114 0 1147 2100
rect 1179 0 1212 2100
rect 1244 0 1277 2100
rect 1309 0 1342 2100
rect 1374 197 1407 2100
rect 4859 1812 5069 1822
rect 4859 1684 5070 1812
rect 4859 1620 4878 1684
rect 4932 1620 5070 1684
rect 4859 1612 5070 1620
rect 4859 1602 5069 1612
rect 1570 1432 4637 1442
rect 1570 1152 1580 1432
rect 1760 1152 2065 1432
rect 2137 1152 2320 1432
rect 2392 1152 2575 1432
rect 2647 1152 2830 1432
rect 2902 1152 3085 1432
rect 3157 1152 3340 1432
rect 3412 1152 4055 1432
rect 4127 1152 4310 1432
rect 4382 1152 4565 1432
rect 4859 1412 5069 1422
rect 4859 1344 5070 1412
rect 4859 1280 4878 1344
rect 4932 1280 5070 1344
rect 4859 1212 5070 1280
rect 4859 1202 5069 1212
rect 1570 1142 4637 1152
rect 4860 1002 5070 1012
rect 2190 992 5070 1002
rect 2190 712 2195 992
rect 2267 712 2453 992
rect 2525 712 2708 992
rect 2780 712 2963 992
rect 3035 712 3218 992
rect 3290 712 3473 992
rect 3545 712 4188 992
rect 4260 712 4443 992
rect 4515 712 4700 992
rect 4752 712 5070 992
rect 2190 702 5070 712
rect 1435 489 1510 497
rect 1435 335 1440 489
rect 1505 335 1510 489
rect 1435 327 1510 335
rect 1840 492 2049 500
rect 1840 292 1848 492
rect 1900 491 2049 492
rect 2041 294 2049 491
rect 3163 482 3247 492
rect 3373 402 3425 412
rect 3478 402 3530 412
rect 3660 402 3740 412
rect 4043 402 4095 412
rect 4148 402 4200 412
rect 4334 404 4440 412
rect 4334 402 4342 404
rect 3247 342 3373 402
rect 3163 332 3373 342
rect 3470 332 3478 402
rect 3530 332 3660 402
rect 3740 332 4043 402
rect 4095 332 4100 402
rect 4145 332 4148 402
rect 4200 340 4342 402
rect 4432 402 4440 404
rect 4728 402 4788 702
rect 4860 692 5070 702
rect 4432 394 4625 402
rect 4432 340 4563 394
rect 4617 340 4625 394
rect 4200 332 4625 340
rect 4678 394 4788 402
rect 4678 340 4686 394
rect 4740 340 4788 394
rect 4678 332 4788 340
rect 4840 492 5070 500
rect 3373 322 3425 332
rect 3478 322 3530 332
rect 3660 322 3740 332
rect 1900 292 2049 294
rect 1840 284 2049 292
rect 4043 285 4095 332
rect 4148 322 4200 332
rect 4840 294 4878 492
rect 5062 294 5070 492
rect 4043 221 4420 285
rect 4840 284 5070 294
rect 1374 187 1458 197
rect 1374 127 1385 187
rect 1449 127 1458 187
rect 1374 117 1458 127
rect 3118 185 3212 194
rect 3118 129 3127 185
rect 3203 129 3212 185
rect 3118 120 3212 129
rect 4355 185 4420 221
rect 4615 185 4685 190
rect 4355 179 4693 185
rect 4355 121 4615 179
rect 4607 120 4615 121
rect 4685 120 4693 179
rect 4607 116 4693 120
<< via2 >>
rect 1580 1152 1760 1432
rect 1443 336 1502 488
rect 1850 297 2038 487
rect 1385 127 1449 187
rect 3127 184 3203 185
rect 3127 130 3128 184
rect 3128 130 3202 184
rect 3202 130 3203 184
rect 3127 129 3203 130
<< metal3 >>
rect 1570 1434 1770 1442
rect 1570 1150 1578 1434
rect 1762 1150 1770 1434
rect 1570 1142 1770 1150
rect 0 489 2048 497
rect 0 335 8 489
rect 292 488 1842 489
rect 292 482 1443 488
rect 292 342 1434 482
rect 292 336 1443 342
rect 1502 336 1842 488
rect 1906 487 2048 489
rect 292 335 1842 336
rect 0 327 1842 335
rect 1840 295 1842 327
rect 2038 297 2048 487
rect 1906 295 2048 297
rect 1840 287 2048 295
rect 1374 189 3017 192
rect 1374 187 2932 189
rect 1374 127 1385 187
rect 1449 127 2932 187
rect 1374 125 2932 127
rect 3009 125 3017 189
rect 1374 122 3017 125
rect 3080 189 3211 196
rect 3080 125 3127 189
rect 3203 125 3211 189
rect 3080 118 3211 125
<< via3 >>
rect 1578 1432 1762 1434
rect 1578 1152 1580 1432
rect 1580 1152 1760 1432
rect 1760 1152 1762 1432
rect 1578 1150 1762 1152
rect 8 335 292 489
rect 1434 342 1443 482
rect 1443 342 1498 482
rect 1842 487 1906 489
rect 1842 297 1850 487
rect 1850 297 1906 487
rect 1842 295 1906 297
rect 2932 125 3009 189
rect 3127 185 3203 189
rect 3127 129 3203 185
rect 3127 125 3203 129
<< metal4 >>
rect 0 497 300 2100
rect 1440 497 1500 2100
rect 0 489 1500 497
rect 0 335 8 489
rect 292 482 1500 489
rect 292 342 1434 482
rect 1498 342 1500 482
rect 292 335 1500 342
rect 0 327 1500 335
rect 0 0 300 327
rect 1440 0 1500 327
rect 1570 1434 1770 2100
rect 1570 1150 1578 1434
rect 1762 1150 1770 1434
rect 1570 0 1770 1150
rect 1840 492 1900 2100
rect 1839 489 1910 492
rect 1839 295 1842 489
rect 1906 295 1910 489
rect 1839 292 1910 295
rect 1840 0 1900 292
rect 2927 189 3208 192
rect 2927 125 2932 189
rect 3009 125 3127 189
rect 3203 125 3208 189
rect 2927 122 3208 125
use sky130_fd_pr__nfet_01v8_9BJ5NV#15tgi  sky130_fd_pr__nfet_01v8_9BJ5NV_1_15tgi
timestamp 1716692466
transform 1 0 4123 0 1 283
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_9BJ5NV#15tgi  sky130_fd_pr__nfet_01v8_9BJ5NV_2_15tgi
timestamp 1716692466
transform 1 0 4651 0 1 281
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_X62NDW#15tgi  sky130_fd_pr__nfet_01v8_lvt_X62NDW_0_15tgi
timestamp 1716692466
transform 1 0 4399 0 1 1072
box -487 -610 487 610
use sky130_fd_pr__pfet_01v8_L75DJ9#15tgi  sky130_fd_pr__pfet_01v8_L75DJ9_0_15tgi
timestamp 1717177055
transform 1 0 3451 0 1 284
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_lvt_E3P74E#15tgi  sky130_fd_pr__pfet_01v8_lvt_E3P74E_0_15tgi
timestamp 1716692466
transform 1 0 2791 0 1 1281
box -871 -819 871 819
<< labels >>
flabel locali 1845 292 2045 492 0 FreeSans 400 0 0 0 VPWR
port 2 nsew power bidirectional
flabel metal2 4870 1612 5070 1812 0 FreeSans 400 0 0 0 EN_N
port 6 nsew signal output
flabel metal2 4870 1212 5070 1412 0 FreeSans 400 0 0 0 EN
port 5 nsew signal output
flabel metal2 4870 292 5070 492 0 FreeSans 400 0 0 0 VGND
port 1 nsew power bidirectional
flabel metal2 4870 702 5070 1002 0 FreeSans 400 0 0 0 AOUT
port 3 nsew analog output
flabel metal2 1570 1142 1770 1442 0 FreeSans 400 0 0 0 AIN
port 4 nsew analog input
flabel metal4 0 327 300 497 0 FreeSans 400 0 0 0 VPWR
port 2 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 5070 2100
<< end >>
